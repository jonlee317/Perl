* File: /net/sim-2/scratch/archive/m_phy/x121/dev/1p0/pyxis/X121/X122_Layout/TOP/X122G001C/X122G001C_CCW.pex.netlist
* Created: Sun Aug 25 10:21:25 2013
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt X122G001C  VDD VSS VSSA_RX VDDHA_RX RXN RXP VDDHA_TX VSSA_TX TXP TXN DO
+ CA0 CA1 CA2 PD PDTX PDRX CCM0 CCM1 CCM2 LBEN DI
* 
XD0_noxref VSS VDD diodenwx  AREA=7.17046e-10 perim=0.00024914 sizedup=0
XD1_noxref VSS VDD diodenwx  AREA=7.17046e-10 perim=0.00024914 sizedup=0
XD2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD10_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD11_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD12_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD13_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD14_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD15_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD16_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD17_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD18_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD19_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD20_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD21_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD22_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD23_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD24_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD25_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD26_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD27_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD28_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD29_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD30_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD31_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD32_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD33_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD34_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD35_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD36_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD37_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD38_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD39_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD40_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD41_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD42_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD43_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD44_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD45_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD46_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD47_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD48_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD49_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD50_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD51_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD52_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD53_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD54_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD55_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD56_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD57_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD58_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD59_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD60_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD61_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD62_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD63_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD64_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD65_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD66_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD67_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD68_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD69_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD70_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD71_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD72_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD73_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD74_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD75_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD76_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD77_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD78_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD79_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD80_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD81_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD82_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD83_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD84_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD85_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD86_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD87_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD88_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD89_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD90_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD91_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD92_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD93_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD94_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD95_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD96_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD97_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD98_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD99_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD100_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD101_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD102_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD103_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD104_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD105_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD106_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD107_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD108_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD109_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD110_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD111_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD112_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD113_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD114_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD115_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD116_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD117_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD118_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XD119_noxref VSS VDD diodenwx  AREA=3.24095e-11 perim=2.332e-05 sizedup=0
XD120_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XD121_noxref VSS VDD diodenwx  AREA=1.32253e-10 perim=5.582e-05 sizedup=0
XD122_noxref VSS VDD diodenwx  AREA=1.32253e-10 perim=5.582e-05 sizedup=0
XD123_noxref VSS VDD diodenwx  AREA=1.32253e-10 perim=5.582e-05 sizedup=0
XD124_noxref VSS VDD diodenwx  AREA=1.32253e-10 perim=5.582e-05 sizedup=0
XD125_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD126_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD127_noxref VSS VDDHA_RX diodenwx  AREA=2.03805e-09 perim=0.00019521 sizedup=0
XD128_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD129_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD130_noxref VSS VDD diodenwx  AREA=4.56213e-10 perim=9.982e-05 sizedup=0
XD131_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD132_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD133_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD134_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD135_noxref VSS VDDHA_RX diodenwx  AREA=2.5624e-09 perim=0.00026291 sizedup=0
XD136_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD137_noxref VSS VDD diodenwx  AREA=4.56213e-10 perim=9.982e-05 sizedup=0
XD138_noxref VSS VDDHA_RX diodenwx  AREA=2.29718e-10 perim=8.804e-05 sizedup=0
XD139_noxref VSS VDD diodenwx  AREA=3.7486e-10 perim=0.00011266 sizedup=0
XD140_noxref VSS VDDHA_RX diodenwx  AREA=3.01127e-10 perim=0.00011624 sizedup=0
XD141_noxref VSS VDDHA_RX diodenwx  AREA=2.29718e-10 perim=8.804e-05 sizedup=0
XD142_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XD143_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782 sizedup=0
XD144_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782 sizedup=0
XD145_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782 sizedup=0
XD146_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782 sizedup=0
XD147_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782 sizedup=0
XD148_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782 sizedup=0
XD149_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782 sizedup=0
XD150_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782 sizedup=0
XD151_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782 sizedup=0
XD152_noxref VSS VDDHA_RX diodenwx  AREA=2.29718e-10 perim=8.804e-05 sizedup=0
XD153_noxref VSS VDD diodenwx  AREA=1.64372e-11 perim=1.641e-05 sizedup=0
XD154_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD155_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD156_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD157_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD158_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD159_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD160_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD161_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD162_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD163_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD164_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD165_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD166_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD167_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD168_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD169_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD170_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD171_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD172_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD173_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD174_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD175_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD176_noxref VSS VDDHA_RX diodenwx  AREA=1.9723e-10 perim=7.73e-05 sizedup=0
XD177_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD178_noxref VSS VDDHA_RX diodenwx  AREA=2.29718e-10 perim=8.804e-05 sizedup=0
XD179_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD180_noxref VSS VDDHA_RX diodenwx  AREA=2.29718e-10 perim=8.804e-05 sizedup=0
XD181_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD182_noxref VSS VDDHA_TX diodenwx  AREA=4.6915e-09 perim=0.00044427 sizedup=0
XD183_noxref VSS VDDHA_RX diodenwx  AREA=2.29718e-10 perim=8.804e-05 sizedup=0
XD184_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD185_noxref VSS VDDHA_RX diodenwx  AREA=2.29718e-10 perim=8.804e-05 sizedup=0
XD186_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XD187_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD188_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD189_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD190_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD191_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD192_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD193_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD194_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD195_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD196_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD197_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD198_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD199_noxref VSS VSSA_TX diodenwx  AREA=2.78358e-09 perim=0.00024351 sizedup=0
XD200_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD201_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD202_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD203_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD204_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD205_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD206_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD207_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD208_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD209_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD210_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD211_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD212_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD213_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD214_noxref VSS VDD diodenwx  AREA=1.64741e-10 perim=6.656e-05 sizedup=0
XD215_noxref VSS VDDHA_TX diodenwx  AREA=2.57441e-08 perim=0.00067856 sizedup=0
XMDC0 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13 PD=1.021e-05
+ PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC0@775 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@774 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@773 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC2 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@121 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@120 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@119 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XX232/D0_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX232/D1_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XMDC0@772 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@771 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@770 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@769 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@768 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@767 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@766 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@765 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@764 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@763 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@762 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@761 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@760 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@759 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@758 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@757 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@756 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@755 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@754 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@753 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@752 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@751 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@750 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@749 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@748 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@747 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@746 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@745 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@744 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@743 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@742 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@741 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@740 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@739 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@738 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@737 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@736 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@735 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@734 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@733 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@732 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@731 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@730 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@729 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@728 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@727 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@726 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@725 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@724 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@723 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@722 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@721 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@720 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@719 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@718 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@717 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@716 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@715 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@714 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@713 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@712 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@711 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@710 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@709 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@708 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@707 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@706 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@705 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@704 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@703 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@702 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@701 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@700 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@699 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@698 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@697 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@696 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@695 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@694 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@693 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@692 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@691 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@690 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@689 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@688 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@687 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@686 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@685 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@684 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@683 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@682 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@681 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@680 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@679 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@678 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@677 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@676 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@675 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@674 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@673 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@672 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@671 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@670 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@669 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@668 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@667 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@666 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@665 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@664 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@663 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@662 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@661 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@660 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@659 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@658 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@657 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@656 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@655 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@654 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@653 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@652 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@651 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@650 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@649 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@648 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@647 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@646 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@645 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@644 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@643 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@642 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@641 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@640 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@639 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@638 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@637 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@636 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@635 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@634 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@633 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@632 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@631 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@630 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@629 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@628 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@627 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@626 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@625 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@624 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@623 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@622 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@621 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@620 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@619 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@618 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@617 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@616 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@615 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@614 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@613 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@612 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@611 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@610 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@609 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@608 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@607 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@606 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@605 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@604 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@603 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@602 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@601 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@600 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@599 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@598 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@597 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@596 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@595 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@594 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@593 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@592 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@591 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@590 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@589 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@588 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@587 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@586 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@585 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@584 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@583 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@582 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@581 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@580 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@579 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@578 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@577 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@576 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@575 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@574 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@573 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@572 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@571 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@570 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@569 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@568 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@567 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@566 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@565 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@564 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@563 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@562 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@561 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@560 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@559 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@558 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@557 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@556 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@555 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@554 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@553 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@552 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@551 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@550 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@549 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@548 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@547 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@546 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@545 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@544 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@543 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@542 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@541 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@540 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@539 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@538 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@537 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@536 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@535 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@534 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@533 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@532 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@531 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@530 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@529 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@528 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@527 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@526 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@525 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@524 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@523 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@522 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@521 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@520 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@519 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@518 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@517 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@516 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@515 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@514 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@513 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@512 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@511 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC2@118 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@117 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@116 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@115 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@114 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@113 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@112 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@111 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@110 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@109 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@108 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@107 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@106 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@105 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@104 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@103 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@102 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@101 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@100 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@99 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@98 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@97 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@96 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@95 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@94 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@93 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@92 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@91 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@90 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@89 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@88 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@87 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@86 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@85 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@84 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@83 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@82 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@81 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@80 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@79 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@78 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@77 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@76 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@75 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@74 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@73 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@72 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@71 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@70 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@69 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@68 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@67 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@66 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@65 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@64 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@63 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@62 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@61 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@60 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@59 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@58 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@57 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@56 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@55 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@54 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@53 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@52 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@51 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@50 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@49 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@48 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@47 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@46 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@45 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@44 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@43 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@42 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@41 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@40 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@39 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@38 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@37 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@36 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@35 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@34 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@33 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@32 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@31 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@30 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@29 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@28 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@27 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@26 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@25 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@24 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@23 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@22 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@21 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@20 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@19 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@18 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XX241/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX241/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX241/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX241/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@510 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@509 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@508 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@507 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@506 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@505 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@504 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@503 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@502 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@501 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@500 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@499 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX242/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX242/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX242/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX242/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@498 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@497 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@496 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@495 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@494 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@493 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX243/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX243/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX243/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX243/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX243/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX243/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX243/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX243/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@492 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@491 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@490 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@489 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@488 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@487 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@486 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@485 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@484 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@483 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@482 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@481 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@480 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@479 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@478 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@477 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@476 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@475 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX244/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX244/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX244/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX244/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX244/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX244/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX244/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX244/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@474 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@473 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@472 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@471 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@470 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@469 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@468 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@467 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@466 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@465 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@464 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@463 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX245/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX245/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX245/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX245/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX245/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX245/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX245/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX245/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@462 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@461 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@460 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@459 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@458 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@457 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@456 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@455 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@454 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@453 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@452 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@451 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX246/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX246/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX246/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX246/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX246/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX246/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX246/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX246/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@450 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@449 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@448 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@447 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@446 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@445 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@444 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@443 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@442 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@441 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@440 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@439 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX247/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX247/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX247/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX247/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX247/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX247/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX247/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX247/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@438 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@437 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@436 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@435 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@434 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@433 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@432 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@431 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@430 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@429 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@428 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@427 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX248/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX248/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX248/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX248/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX248/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX248/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX248/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX248/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@426 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@425 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@424 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@423 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@422 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@421 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@420 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@419 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@418 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@417 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@416 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@415 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX249/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX249/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX249/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX249/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX249/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX249/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX249/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX249/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@414 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@413 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@412 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@411 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@410 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@409 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@408 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@407 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@406 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@405 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@404 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@403 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX250/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX250/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX250/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX250/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX250/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX250/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX250/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX250/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@402 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@401 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@400 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@399 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@398 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@397 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@396 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@395 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@394 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@393 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@392 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@391 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX251/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX251/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX251/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX251/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX251/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX251/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX251/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX251/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@390 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@389 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@388 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@387 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@386 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@385 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@384 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@383 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@382 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@381 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@380 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@379 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX252/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX252/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX252/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX252/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX252/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX252/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX252/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX252/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@378 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@377 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@376 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@375 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@374 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@373 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@372 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@371 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@370 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@369 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@368 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@367 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX253/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX253/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX253/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX253/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX253/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX253/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX253/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX253/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@366 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@365 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@364 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@363 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@362 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@361 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@360 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@359 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@358 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@357 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@356 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@355 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX254/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D10_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D11_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D12_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D13_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D14_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX254/D15_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@354 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@353 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@352 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@351 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@350 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@349 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@348 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@347 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@346 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@345 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@344 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@343 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@342 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@341 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@340 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@339 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@338 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@337 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@336 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@335 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@334 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@333 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@332 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@331 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX255/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX255/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX255/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX255/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@330 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@329 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@328 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@327 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@326 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@325 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX256/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX256/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX256/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX256/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX256/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@324 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@323 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@322 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@321 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@320 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@319 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@318 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@317 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@316 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@315 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX257/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX257/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX257/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX257/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX257/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@314 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@313 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@312 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@311 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@310 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX258/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX258/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX258/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX258/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX258/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX258/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX258/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX258/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX258/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX258/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@309 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@308 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@307 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@306 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@305 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@304 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@303 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@302 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@301 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@300 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@299 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@298 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@297 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@296 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@295 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX259/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX259/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX259/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX259/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX259/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX259/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX259/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX259/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX259/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX259/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@294 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@293 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@292 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@291 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@290 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@289 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@288 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@287 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@286 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@285 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX260/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX260/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX260/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX260/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX260/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX260/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX260/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX260/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX260/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX260/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@284 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@283 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@282 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@281 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@280 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@279 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@278 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@277 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@276 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@275 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX261/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX261/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX261/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX261/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX261/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX261/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX261/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX261/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX261/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX261/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@274 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@273 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@272 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@271 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@270 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@269 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@268 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@267 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@266 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@265 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX262/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX262/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX262/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX262/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX262/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX262/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX262/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX262/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX262/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX262/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@264 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@263 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@262 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@261 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@260 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@259 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@258 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@257 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@256 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@255 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX263/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX263/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX263/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX263/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX263/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX263/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX263/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX263/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX263/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX263/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@254 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@253 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@252 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@251 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@250 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@249 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@248 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@247 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@246 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@245 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX264/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX264/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX264/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX264/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX264/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX264/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX264/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX264/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX264/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX264/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@244 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@243 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@242 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@241 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@240 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@239 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@238 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@237 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@236 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@235 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX265/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX265/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX265/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX265/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX265/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX265/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX265/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX265/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX265/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX265/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@234 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@233 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@232 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@231 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@230 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@229 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@228 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@227 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@226 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@225 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX266/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX266/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX266/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX266/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX266/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX266/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX266/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX266/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX266/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX266/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@224 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@223 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@222 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@221 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@220 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@219 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@218 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@217 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@216 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@215 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX267/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX267/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX267/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX267/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX267/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX267/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX267/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX267/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX267/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX267/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@214 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@213 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@212 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@211 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@210 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@209 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@208 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@207 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@206 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@205 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX268/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX268/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX268/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX268/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX268/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX268/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX268/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX268/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX268/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX268/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@204 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@203 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@202 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@201 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@200 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@199 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@198 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@197 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@196 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@195 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX269/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D5_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D6_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D7_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D8_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D9_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D10_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D11_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D12_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D13_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D14_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D15_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D16_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D17_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D18_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX269/D19_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@194 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@193 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@192 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@191 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@190 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@189 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@188 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@187 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@186 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@185 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@184 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@183 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@182 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@181 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@180 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@179 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@178 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@177 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@176 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@175 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX270/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX270/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX270/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX270/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX270/D4_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@174 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@173 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@172 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@171 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@170 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX271/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@169 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@168 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@167 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@166 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX272/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@165 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@164 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX273/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX273/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@163 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@162 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@161 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@160 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@159 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@158 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX274/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX274/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@157 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@156 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@155 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@154 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX275/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX275/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@153 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@152 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@151 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@150 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX276/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX276/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@149 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@148 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@147 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@146 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX277/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX277/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@145 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@144 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@143 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@142 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX278/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX278/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@141 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@140 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@139 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@138 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@137 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@136 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@135 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@134 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX279/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@133 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@132 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@131 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@130 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@129 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@128 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@127 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@126 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX280/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX280/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@125 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@124 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@123 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@122 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@121 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@120 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@119 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@118 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@117 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@116 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@115 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@114 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@113 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@112 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@111 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@110 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@109 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@108 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX282/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX282/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@107 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@106 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@105 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@104 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@103 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@102 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@101 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@100 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@99 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@98 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX283/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX283/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@97 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@96 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@95 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@94 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@93 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@92 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@91 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@90 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX284/D0_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX284/D1_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX284/D2_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XX284/D3_noxref VSS VDD diodenwx  AREA=3.47875e-11 perim=2.36e-05 sizedup=0
XMDC0@89 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@88 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@87 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@86 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@85 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@84 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@83 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@82 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@81 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@80 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@79 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@78 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@77 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@76 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@75 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@74 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@73 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@72 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@71 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@70 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@69 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@68 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=10.511 scb=0.0093744 scc=0.000692813
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX286/D0_noxref VDDHA_RX VDDHA_RX egdiodepnw  AREA=2.496e-13 perim=6.4e-06
+ sizedup=0
XX286/D1_noxref VDDHA_RX VDDHA_RX egdiodepnw  AREA=4.088e-13 perim=1.038e-05
+ sizedup=0
XX286/D2_noxref VDDHA_RX VDDHA_RX egdiodepnw  AREA=4.088e-13 perim=1.038e-05
+ sizedup=0
XX286/D3_noxref VDDHA_RX VDDHA_RX egdiodepnw  AREA=4.088e-13 perim=1.038e-05
+ sizedup=0
XX286/D4_noxref VDDHA_RX VDDHA_RX egdiodepnw  AREA=4.088e-13 perim=1.038e-05
+ sizedup=0
XX286/D5_noxref VSS VDD diodenwx  AREA=4.51385e-12 perim=8.85e-06 sizedup=0
XX286/D6_noxref VSS VDDHA_RX diodenwx  AREA=8.24875e-11 perim=3.643e-05
+ sizedup=0
XX286/D7_noxref VSS VDD diodenwx  AREA=1.4999e-11 perim=1.562e-05 sizedup=0
XX286/D8_noxref VSS VDDHA_RX diodenwx  AREA=2.61907e-10 perim=9.677e-05
+ sizedup=0
XX286/D9_noxref VSS VDDHA_RX diodenwx  AREA=4.47156e-10 perim=0.00012697
+ sizedup=0
XX286/D10_noxref VSS VDD diodenwx  AREA=3.00641e-11 perim=2.246e-05 sizedup=0
XX286/D11_noxref VSS VDDHA_RX diodenwx  AREA=7.4885e-11 perim=4.281e-05
+ sizedup=0
XX286/D12_noxref VSS VDD diodenwx  AREA=5.15602e-11 perim=3.169e-05 sizedup=0
XX286/D13_noxref VSS VDDHA_RX diodenwx  AREA=1.66066e-10 perim=5.382e-05
+ sizedup=0
XX286/D14_noxref VSS VDDHA_RX diodenwx  AREA=3.11259e-10 perim=8.664e-05
+ sizedup=0
XX286/D15_noxref VSS VDDHA_RX diodenwx  AREA=2.61907e-10 perim=9.677e-05
+ sizedup=0
XX286/D16_noxref VSS VDDHA_RX diodenwx  AREA=1.83562e-10 perim=5.708e-05
+ sizedup=0
XXI1/XI3/XG3B/M4 XI1/XI3/XG3B/N1 XI1/XI3/TIEL VSS VSS nfet L=3e-08 W=1.26e-06
+ AD=7.56e-14 AS=1.323e-13 PD=1.38e-06 PS=2.73e-06 M=1 sca=2.20935
+ scb=0.000220603 scc=4.87494e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06
+ sa=1.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG3B/M3 XI1/XI3/N3B XI1/XI3/N2B XI1/XI3/XG3B/N1 VSS nfet L=3e-08
+ W=1.26e-06 AD=1.323e-13 AS=7.56e-14 PD=2.73e-06 PS=1.38e-06 M=1 sca=2.02283
+ scb=0.000138581 scc=1.6485e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06
+ sa=2.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG6B/M2 XI1/XI3/N2A XI1/XI3/N2B VSS VSS nfet L=3e-08 W=3.2e-07
+ AD=3.36e-14 AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=1.04999 scb=5.83778e-05
+ scc=3.95488e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG2B/M2 XI1/XI3/N2B XI1/XI3/N1B VSS VSS nfet L=3e-08 W=3.2e-07
+ AD=3.36e-14 AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=1.04999 scb=5.83778e-05
+ scc=3.95488e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG5B/M2 XI1/XI3/N1A XI1/XI3/N1B VSS VSS nfet L=3e-08 W=3.2e-07
+ AD=3.36e-14 AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=1.04999 scb=5.83778e-05
+ scc=3.95488e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG1B/M2 XI1/XI3/N1B XI1/NN VSS VSS nfet L=3e-08 W=3.2e-07 AD=3.36e-14
+ AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=1.04999 scb=5.83778e-05
+ scc=3.95488e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG1A/M2 XI1/XI3/N1A XI1/NP VSS VSS nfet L=3e-08 W=3.2e-07 AD=3.36e-14
+ AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=1.04999 scb=5.83778e-05
+ scc=3.95488e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG5A/M2 XI1/XI3/N1B XI1/XI3/N1A VSS VSS nfet L=3e-08 W=3.2e-07
+ AD=3.36e-14 AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=1.04999 scb=5.83778e-05
+ scc=3.95488e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG2A/M2 XI1/XI3/N2A XI1/XI3/N1A VSS VSS nfet L=3e-08 W=3.2e-07
+ AD=3.36e-14 AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=1.04999 scb=5.83778e-05
+ scc=3.95488e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG6A/M2 XI1/XI3/N2B XI1/XI3/N2A VSS VSS nfet L=3e-08 W=3.2e-07
+ AD=3.36e-14 AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=1.04999 scb=5.83778e-05
+ scc=3.95488e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG3A/M3 XI1/XI3/N3A XI1/XI3/N2A XI1/XI3/XG3A/N1 VSS nfet L=3e-08
+ W=1.26e-06 AD=1.323e-13 AS=7.56e-14 PD=2.73e-06 PS=1.38e-06 M=1 sca=0.771574
+ scb=2.1376e-05 scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06
+ sa=1.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG3A/M4 XI1/XI3/XG3A/N1 XI1/VAL VSS VSS nfet L=3e-08 W=1.26e-06
+ AD=7.56e-14 AS=1.323e-13 PD=1.38e-06 PS=2.73e-06 M=1 sca=0.771574
+ scb=2.1376e-05 scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06
+ sa=2.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XMDC2@17 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@16 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG3B/M2 XI1/XI3/N3B XI1/XI3/TIEL VDD VDD pfet L=3e-08 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=31.4978 scb=0.0263811
+ scc=0.0031947 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=2.55e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI3/XG3B/M1 XI1/XI3/N3B XI1/XI3/N2B VDD VDD pfet L=3e-08 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=30.0289 scb=0.0235667
+ scc=0.00309381 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=2.55e-07 sb=1.05e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI3/XG6B/M1 XI1/XI3/N2A XI1/XI3/N2B VDD VDD pfet L=3e-08 W=9.6e-07
+ AD=1.008e-13 AS=1.008e-13 PD=2.13e-06 PS=2.13e-06 M=1 sca=29.0612
+ scb=0.0206647 scc=0.0031671 lpccnr=3.1e-08 covpccnr=0 wrxcnr=8.64e-07
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG2B/M1 XI1/XI3/N2B XI1/XI3/N1B VDD VDD pfet L=3e-08 W=9.6e-07
+ AD=1.008e-13 AS=1.008e-13 PD=2.13e-06 PS=2.13e-06 M=1 sca=29.4128
+ scb=0.0213427 scc=0.00317186 lpccnr=3.1e-08 covpccnr=0 wrxcnr=8.64e-07
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG5B/M1 XI1/XI3/N1A XI1/XI3/N1B VDD VDD pfet L=3e-08 W=3.2e-07
+ AD=3.36e-14 AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=62.7891 scb=0.0436616
+ scc=0.00843965 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG1B/M1 XI1/XI3/N1B XI1/NN VDD VDD pfet L=3e-08 W=3.2e-07 AD=3.36e-14
+ AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=75.786 scb=0.0575399 scc=0.0109618
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI3/XG1A/M1 XI1/XI3/N1A XI1/NP VDD VDD pfet L=3e-08 W=3.2e-07 AD=3.36e-14
+ AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=75.786 scb=0.0575399 scc=0.0109618
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI3/XG5A/M1 XI1/XI3/N1B XI1/XI3/N1A VDD VDD pfet L=3e-08 W=3.2e-07
+ AD=3.36e-14 AS=3.36e-14 PD=8.5e-07 PS=8.5e-07 M=1 sca=62.7891 scb=0.0436616
+ scc=0.00843965 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.88e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG2A/M1 XI1/XI3/N2A XI1/XI3/N1A VDD VDD pfet L=3e-08 W=9.6e-07
+ AD=1.008e-13 AS=1.008e-13 PD=2.13e-06 PS=2.13e-06 M=1 sca=27.8184
+ scb=0.0210548 scc=0.00317176 lpccnr=3.1e-08 covpccnr=0 wrxcnr=8.64e-07
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG6A/M1 XI1/XI3/N2B XI1/XI3/N2A VDD VDD pfet L=3e-08 W=9.6e-07
+ AD=1.008e-13 AS=1.008e-13 PD=2.13e-06 PS=2.13e-06 M=1 sca=26.7929
+ scb=0.0197965 scc=0.00316597 lpccnr=3.1e-08 covpccnr=0 wrxcnr=8.64e-07
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG3A/M1 XI1/XI3/N3A XI1/XI3/N2A VDD VDD pfet L=3e-08 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=25.1334 scb=0.0186433
+ scc=0.00304011 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=2.55e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI3/XG3A/M2 XI1/XI3/N3A XI1/VAL VDD VDD pfet L=3e-08 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=24.9886 scb=0.0186011
+ scc=0.0030401 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=2.55e-07 sb=1.05e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC1 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=5.56363 scb=0.00460522
+ scc=0.000177115 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@2 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@3 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@4 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@5 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@6 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@7 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=5.54632 scb=0.00458332
+ scc=0.000175109 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC0 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06
+ PS=1.024e-05 M=1 sca=2.17718 scb=0.00103367 scc=1.0163e-05 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC0@28 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/MDC1@8 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=5.54632 scb=0.00458332
+ scc=0.000175109 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC0@27 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/MDC1@9 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC0@26 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/MDC1@10 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC0@25 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/MDC1@11 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC0@24 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/MDC1@12 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC0@23 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=6e-13 AS=3.5e-13
+ PD=1.024e-05 PS=5.14e-06 M=1 sca=2.17718 scb=0.00103367 scc=1.0163e-05
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/MDC1@13 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@14 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6862 scb=0.00304112
+ scc=0.000115443 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@15 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=5.56363 scb=0.00460522
+ scc=0.000177115 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/RRP XI1/INPI RXP VDDHA_RX opppcres 231.017 M=1 w=2.945e-06 l=1e-06 bp=1
+ pbar=1 s=1 ncr=1 sizedup=0 
XXI1/M2P XI1/INPI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06 AD=1.75e-13
+ AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1 sca=0.995619 scb=0.000146103
+ scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M2P@8 XI1/INPI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=6.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2P@7 XI1/INPI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=1.1e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2P@6 XI1/INPI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=1.59e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2P@5 XI1/INPI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=2.0083e-06 sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2P@4 XI1/INPI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=2.0083e-06 sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2P@3 XI1/INPI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=2.0083e-06 sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2P@2 XI1/INPI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1 sca=0.995619 scb=0.000146103
+ scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1P XI1/INPI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1 sca=12.0388 scb=0.0126667
+ scc=0.000383588 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1P@8 XI1/INPI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=7.16658 scb=0.00451039
+ scc=3.53414e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=6.1e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1P@7 XI1/INPI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=5.63416 scb=0.0026305
+ scc=2.42385e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=1.1e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1P@6 XI1/INPI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=4.95944 scb=0.00226274
+ scc=2.3935e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=1.59e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1P@5 XI1/INPI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=3.83107 scb=0.00218279
+ scc=2.39272e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=2.0083e-06
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1P@4 XI1/INPI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=3.83107 scb=0.00218279
+ scc=2.39272e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=2.0083e-06
+ sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1P@3 XI1/INPI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=3.83107 scb=0.00218279
+ scc=2.39272e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=2.0083e-06
+ sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1P@2 XI1/INPI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1 sca=3.83107 scb=0.00218279
+ scc=2.39272e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/RRN XI1/INNI RXN VDDHA_RX opppcres 231.017 M=1 w=2.945e-06 l=1e-06   bp=1
+ pbar=1 s=1 ncr=1 sizedup=0
XXI1/M2N XI1/INNI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06 AD=1.75e-13
+ AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1 sca=0.995619 scb=0.000146103
+ scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M2N@8 XI1/INNI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=6.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2N@7 XI1/INNI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=1.1e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2N@6 XI1/INNI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=1.59e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2N@5 XI1/INNI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=2.0083e-06 sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2N@4 XI1/INNI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=2.0083e-06 sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2N@3 XI1/INNI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=0.995619
+ scb=0.000146103 scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06
+ sa=2.0083e-06 sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/M2N@2 XI1/INNI VSSA_RX VSSA_RX VSSA_RX egnfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1 sca=0.995619 scb=0.000146103
+ scc=1.37973e-07 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1N XI1/INNI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1 sca=12.0388 scb=0.0126667
+ scc=0.000383588 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1N@8 XI1/INNI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=7.16658 scb=0.00451039
+ scc=3.53414e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=6.1e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1N@7 XI1/INNI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=5.63416 scb=0.0026305
+ scc=2.42385e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=1.1e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1N@6 XI1/INNI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=4.95944 scb=0.00226274
+ scc=2.3935e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=1.59e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1N@5 XI1/INNI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=3.83107 scb=0.00218279
+ scc=2.39272e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=2.0083e-06
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1N@4 XI1/INNI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=3.83107 scb=0.00218279
+ scc=2.39272e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=2.0083e-06
+ sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1N@3 XI1/INNI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=3.83107 scb=0.00218279
+ scc=2.39272e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=2.0083e-06
+ sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/M1N@2 XI1/INNI VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.5e-06
+ AD=1.75e-13 AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1 sca=3.83107 scb=0.00218279
+ scc=2.39272e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.25e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M3N XI1/XI1/N2N XI1/XI1/N1P VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.05e-07
+ sb=2.0022e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M3N@4 XI1/XI1/N2N XI1/XI1/N1P VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=4.75e-07
+ sb=2.0022e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M3N@3 XI1/XI1/N2N XI1/XI1/N1P VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=8.45e-07
+ sb=1.955e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M3N@2 XI1/XI1/N2N XI1/XI1/N1P VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.215e-06
+ sb=1.585e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M2N XI1/XI1/N1P XI1/XI1/N1P VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.585e-06
+ sb=1.215e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M2N@4 XI1/XI1/N1P XI1/XI1/N1P VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.955e-06
+ sb=8.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M2N@3 XI1/XI1/N1P XI1/XI1/N1P VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0022e-06
+ sb=4.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M2N@2 XI1/XI1/N1P XI1/XI1/N1P VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0022e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M12N XI1/XI1/N1P XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0.90884 scb=3.09084e-05
+ scc=1.0981e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI1/M4N XI1/XI1/N2N XI1/XI1/N2N VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=7.0669
+ scb=0.00557941 scc=0.000311232 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.05e-07 sb=1.995e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M4N@4 XI1/XI1/N2N XI1/XI1/N2N VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=3.75e-07 sb=1.725e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M4N@3 XI1/XI1/N2N XI1/XI1/N2N VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=6.45e-07 sb=1.455e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M4N@2 XI1/XI1/N2N XI1/XI1/N2N VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=9.15e-07 sb=1.185e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M5N XI1/INP1 XI1/XI1/N2N VDD VDD pfet L=1.5e-07 W=3.54e-06 AD=2.124e-13
+ AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386 scb=0.00553092
+ scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06 sa=1.185e-06
+ sb=9.15e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M5N@4 XI1/INP1 XI1/XI1/N2N VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.455e-06 sb=6.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M5N@3 XI1/INP1 XI1/XI1/N2N VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.725e-06 sb=3.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M5N@2 XI1/INP1 XI1/XI1/N2N VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.995e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M0 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@24 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=5.4e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@23 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=9.6e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M11N XI1/XI1/N2N XI1/XI1/PDB VDD VDD egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=24.4822 scb=0.0304636
+ scc=0.00212873 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI1/M1N XI1/XI1/N1P XI1/INNI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@22 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=1.38e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1N@8 XI1/XI1/N1P XI1/INNI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=5.6e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@21 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=1.8e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1N@7 XI1/XI1/N1P XI1/INNI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@20 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@19 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1N@6 XI1/XI1/N1P XI1/INNI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.44e-06
+ sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@18 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=1.8e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1N@5 XI1/XI1/N1P XI1/INNI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.88e-06
+ sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@17 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=1.38e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1N@4 XI1/XI1/N1P XI1/INNI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI1/M0@16 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=9.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1N@3 XI1/XI1/N1P XI1/INNI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@15 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1N@2 XI1/XI1/N1P XI1/INNI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@14 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M7P XI1/INP1 XI1/INN1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=1.645e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M7P@4 XI1/INP1 XI1/INN1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=3.25e-07 sb=1.425e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M7P@3 XI1/INP1 XI1/INN1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=5.45e-07 sb=1.205e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M7P@2 XI1/INP1 XI1/INN1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=7.65e-07 sb=9.85e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M6N XI1/INP1 XI1/INP1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=9.85e-07 sb=7.65e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M6N@4 XI1/INP1 XI1/INP1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.205e-06 sb=5.45e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M6N@3 XI1/INP1 XI1/INP1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.425e-06 sb=3.25e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M6N@2 XI1/INP1 XI1/INP1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.645e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M10N XI1/INP1 XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M3P XI1/XI1/N2P XI1/XI1/N1N VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.05e-07
+ sb=2.0022e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M3P@4 XI1/XI1/N2P XI1/XI1/N1N VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=4.75e-07
+ sb=2.0022e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M3P@3 XI1/XI1/N2P XI1/XI1/N1N VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=8.45e-07
+ sb=1.955e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M3P@2 XI1/XI1/N2P XI1/XI1/N1N VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.215e-06
+ sb=1.585e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M2P XI1/XI1/N1N XI1/XI1/N1N VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.585e-06
+ sb=1.215e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M2P@4 XI1/XI1/N1N XI1/XI1/N1N VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.955e-06
+ sb=8.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M2P@3 XI1/XI1/N1N XI1/XI1/N1N VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0022e-06
+ sb=4.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M2P@2 XI1/XI1/N1N XI1/XI1/N1N VSSA_RX VSSA_RX nfet L=2.5e-07 W=4e-06
+ AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1 sca=1.23045 scb=0.000159171
+ scc=2.70528e-07 lpccnr=2.29e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0022e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/X1I291/M2 XI1/XI1/PDB XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M12P XI1/XI1/N1N XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0.90884 scb=3.09084e-05
+ scc=1.0981e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI1/M4P XI1/XI1/N2P XI1/XI1/N2P VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=7.0669
+ scb=0.00557941 scc=0.000311232 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.05e-07 sb=1.995e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M4P@4 XI1/XI1/N2P XI1/XI1/N2P VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=3.75e-07 sb=1.725e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M4P@3 XI1/XI1/N2P XI1/XI1/N2P VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=6.45e-07 sb=1.455e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M4P@2 XI1/XI1/N2P XI1/XI1/N2P VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=9.15e-07 sb=1.185e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M5P XI1/INN1 XI1/XI1/N2P VDD VDD pfet L=1.5e-07 W=3.54e-06 AD=2.124e-13
+ AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386 scb=0.00553092
+ scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06 sa=1.185e-06
+ sb=9.15e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M5P@4 XI1/INN1 XI1/XI1/N2P VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.455e-06 sb=6.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M5P@3 XI1/INN1 XI1/XI1/N2P VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.725e-06 sb=3.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M5P@2 XI1/INN1 XI1/XI1/N2P VDD VDD pfet L=1.5e-07 W=3.54e-06
+ AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=6.05386
+ scb=0.00553092 scc=0.000311229 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.995e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/X1I291/M1 XI1/XI1/PDB XI1/PDI VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=5.76429
+ scb=0.00422298 scc=3.53586e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M0@13 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@12 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=5.4e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@11 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=9.6e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M11P XI1/XI1/N2P XI1/XI1/PDB VDD VDD egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=24.4822 scb=0.0304636
+ scc=0.00212873 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI1/M1P XI1/XI1/N1N XI1/INPI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@10 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=1.38e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1P@8 XI1/XI1/N1N XI1/INPI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=5.6e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@9 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=1.8e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1P@7 XI1/XI1/N1N XI1/INPI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@8 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@7 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1P@6 XI1/XI1/N1N XI1/INPI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.44e-06
+ sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@6 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=1.8e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1P@5 XI1/XI1/N1N XI1/INPI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.88e-06
+ sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@5 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=1.38e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1P@4 XI1/XI1/N1N XI1/INPI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI1/M0@4 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=9.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1P@3 XI1/XI1/N1N XI1/INPI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@3 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M1P@2 XI1/XI1/N1N XI1/INPI XI1/XI1/N0 VDDHA_RX egpfet L=3e-07 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.9497 scb=0.00165427
+ scc=7.03629e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M0@2 XI1/XI1/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=3.33827 scb=0.00278801
+ scc=5.32744e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI1/M7N XI1/INN1 XI1/INP1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=1.645e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M7N@4 XI1/INN1 XI1/INP1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=3.25e-07 sb=1.425e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M7N@3 XI1/INN1 XI1/INP1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=5.45e-07 sb=1.205e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M7N@2 XI1/INN1 XI1/INP1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=7.65e-07 sb=9.85e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M6P XI1/INN1 XI1/INN1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=9.85e-07 sb=7.65e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M6P@4 XI1/INN1 XI1/INN1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.205e-06 sb=5.45e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M6P@3 XI1/INN1 XI1/INN1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.425e-06 sb=3.25e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M6P@2 XI1/INN1 XI1/INN1 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.645e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI1/M10P XI1/INN1 XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M3P XI1/XI5/XI0B/N2P XI1/XI5/XI0B/N1N VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.05e-07 sb=1.215e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M3P@2 XI1/XI5/XI0B/N2P XI1/XI5/XI0B/N1N VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=4.75e-07 sb=8.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M2P XI1/XI5/XI0B/N1N XI1/XI5/XI0B/N1N VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=8.45e-07 sb=4.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M2P@2 XI1/XI5/XI0B/N1N XI1/XI5/XI0B/N1N VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.215e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M2N XI1/XI5/XI0B/N1P XI1/XI5/XI0B/N1P VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.05e-07 sb=1.215e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M2N@2 XI1/XI5/XI0B/N1P XI1/XI5/XI0B/N1P VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=4.75e-07 sb=8.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M3N XI1/XI5/XI0B/N2N XI1/XI5/XI0B/N1P VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=8.45e-07 sb=4.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M3N@2 XI1/XI5/XI0B/N2N XI1/XI5/XI0B/N1P VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.215e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XX286/X72/X8/D0_noxref VSS VDD diodenwx  AREA=4.11324e-11 perim=2.72e-05
+ sizedup=0
XXI1/XI5/XI0B/M5P XI1/XI5/XI0B/N3N XI1/XI5/XI0B/N2P VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=7.53851
+ scb=0.00589959 scc=0.000336008 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.05e-07 sb=9.15e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M5P@2 XI1/XI5/XI0B/N3N XI1/XI5/XI0B/N2P VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=7.27107
+ scb=0.00581659 scc=0.00033599 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=3.75e-07 sb=6.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M4P XI1/XI5/XI0B/N2P XI1/XI5/XI0B/N2P VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.24568
+ scb=0.0057654 scc=0.000335987 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=6.45e-07 sb=3.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M4P@2 XI1/XI5/XI0B/N2P XI1/XI5/XI0B/N2P VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=6.24568
+ scb=0.0057654 scc=0.000335987 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=9.15e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M14P XI1/XI5/XI0B/N1N422 XI1/XI5/XI0B/N1N422 VDD VDD pfet
+ L=1.8e-07 W=2e-06 AD=1.2e-13 AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1
+ sca=3.38053 scb=0.00159701 scc=1.61519e-05 lpccnr=1.66e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.05e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M14P@2 XI1/XI5/XI0B/N1N422 XI1/XI5/XI0B/N1N422 VDD VDD pfet
+ L=1.8e-07 W=2e-06 AD=1.2e-13 AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1
+ sca=3.38053 scb=0.00159701 scc=1.61519e-05 lpccnr=1.66e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M14N XI1/XI5/O2 XI1/XI5/XI0B/N1N422 VDD VDD pfet L=1.8e-07 W=2e-06
+ AD=1.2e-13 AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1 sca=3.38053 scb=0.00159701
+ scc=1.61519e-05 lpccnr=1.66e-07 covpccnr=0 wrxcnr=1.8e-06 sa=1.05e-07
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M14N@2 XI1/XI5/O2 XI1/XI5/XI0B/N1N422 VDD VDD pfet L=1.8e-07
+ W=2e-06 AD=1.2e-13 AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1 sca=3.38053
+ scb=0.00159701 scc=1.61519e-05 lpccnr=1.66e-07 covpccnr=0 wrxcnr=1.8e-06
+ sa=4.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M4N XI1/XI5/XI0B/N2N XI1/XI5/XI0B/N2N VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=6.24568
+ scb=0.0057654 scc=0.000335987 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.05e-07 sb=9.15e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M4N@2 XI1/XI5/XI0B/N2N XI1/XI5/XI0B/N2N VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.24568
+ scb=0.0057654 scc=0.000335987 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=3.75e-07 sb=6.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M5N XI1/XI5/XI0B/N3P XI1/XI5/XI0B/N2N VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=7.27107
+ scb=0.00581659 scc=0.00033599 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=6.45e-07 sb=3.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M5N@2 XI1/XI5/XI0B/N3P XI1/XI5/XI0B/N2N VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=7.53851
+ scb=0.00589959 scc=0.000336008 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=9.15e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/MDC3 VDDHA_RX IBRX2 VDDHA_RX VDDHA_RX egpfet L=2e-06 W=6e-06
+ AD=7.2e-13 AS=7.2e-13 PD=1.224e-05 PS=1.224e-05 M=1 sca=4 scb=0.00306566
+ scc=0.000422923 lpccnr=1.815e-06 covpccnr=0 wrxcnr=5.4e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/X1I291/M1 XI1/XI5/XI0B/PDB XI1/PDI VDDHA_RX VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=1.70503 scb=0.000376785 scc=2.23221e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M11P XI1/XI5/XI0B/N2P XI1/XI5/XI0B/PDB VDD VDD egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=18.5703
+ scb=0.0243185 scc=0.000992376 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M1I437 XI1/XI5/XI0B/N1N422 XI1/XI5/XI0B/PDB VDD VDD egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=16.5926 scb=0.0212421 scc=0.000750386 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M1P XI1/XI5/XI0B/N1N IBRX2 XI1/XI5/XI0B/N0 VDDHA_RX egpfet L=3e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0@12 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=5.4e-07 sb=1.8e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0@11 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=9.6e-07 sb=1.38e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M1P@4 XI1/XI5/XI0B/N1N IBRX2 XI1/XI5/XI0B/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=5.6e-07 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0@10 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.38e-06 sb=9.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M1P@3 XI1/XI5/XI0B/N1N IBRX2 XI1/XI5/XI0B/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0@9 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.8e-06 sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M1P@2 XI1/XI5/XI0B/N1N IBRX2 XI1/XI5/XI0B/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.44e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0@8 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0@7 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M1N XI1/XI5/XI0B/N1P XI1/INNI XI1/XI5/XI0B/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0@6 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=5.4e-07 sb=1.8e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M1N@4 XI1/XI5/XI0B/N1P XI1/INNI XI1/XI5/XI0B/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=5.6e-07 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0@5 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=9.6e-07 sb=1.38e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0@4 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.38e-06 sb=9.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M1N@3 XI1/XI5/XI0B/N1P XI1/INNI XI1/XI5/XI0B/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0@3 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.8e-06 sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M1N@2 XI1/XI5/XI0B/N1P XI1/INNI XI1/XI5/XI0B/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.44e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M0@2 XI1/XI5/XI0B/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M11N XI1/XI5/XI0B/N2N XI1/XI5/XI0B/PDB VDD VDD egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=18.5703
+ scb=0.0243185 scc=0.000992376 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M7N XI1/XI5/XI0B/N3N XI1/XI5/XI0B/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=1.005e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0B/M7N@2 XI1/XI5/XI0B/N3N XI1/XI5/XI0B/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=4.05e-07 sb=7.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0B/M6P XI1/XI5/XI0B/N3N XI1/XI5/XI0B/N3N VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=7.05e-07 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0B/M6P@2 XI1/XI5/XI0B/N3N XI1/XI5/XI0B/N3N VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.005e-06 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0B/M13P XI1/XI5/XI0B/N1N422 XI1/XI5/XI0B/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0B/M13P@2 XI1/XI5/XI0B/N1N422 XI1/XI5/XI0B/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=4.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0B/M10P XI1/XI5/XI0B/N3N XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M12P XI1/XI5/XI0B/N1N XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M7P XI1/XI5/XI0B/N3P XI1/XI5/XI0B/N3N VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=1.005e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0B/M7P@2 XI1/XI5/XI0B/N3P XI1/XI5/XI0B/N3N VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=4.05e-07 sb=7.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0B/M6N XI1/XI5/XI0B/N3P XI1/XI5/XI0B/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=7.05e-07 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0B/M6N@2 XI1/XI5/XI0B/N3P XI1/XI5/XI0B/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.005e-06 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0B/M13N XI1/XI5/O2 XI1/XI5/XI0B/N3N VSSA_RX VSSA_RX nfet L=1.8e-07
+ W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=4.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M13N@2 XI1/XI5/O2 XI1/XI5/XI0B/N3N VSSA_RX VSSA_RX nfet L=1.8e-07
+ W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=4.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M10N XI1/XI5/XI0B/N3P XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/M12N XI1/XI5/XI0B/N1P XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/X1I291/M2 XI1/XI5/XI0B/PDB XI1/PDI VSSA_RX VSSA_RX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0B/M13 XI1/XI5/O2 XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M3P XI1/XI5/XI0A/N2P XI1/XI5/XI0A/N1N VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.05e-07 sb=1.215e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M3P@2 XI1/XI5/XI0A/N2P XI1/XI5/XI0A/N1N VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=4.75e-07 sb=8.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M2P XI1/XI5/XI0A/N1N XI1/XI5/XI0A/N1N VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=8.45e-07 sb=4.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M2P@2 XI1/XI5/XI0A/N1N XI1/XI5/XI0A/N1N VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.215e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M2N XI1/XI5/XI0A/N1P XI1/XI5/XI0A/N1P VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.05e-07 sb=1.215e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M2N@2 XI1/XI5/XI0A/N1P XI1/XI5/XI0A/N1P VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=4.75e-07 sb=8.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M3N XI1/XI5/XI0A/N2N XI1/XI5/XI0A/N1P VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=2.4e-13 PD=4.12e-06 PS=4.12e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=8.45e-07 sb=4.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M3N@2 XI1/XI5/XI0A/N2N XI1/XI5/XI0A/N1P VSSA_RX VSSA_RX nfet
+ L=2.5e-07 W=4e-06 AD=2.4e-13 AS=4.2e-13 PD=4.12e-06 PS=8.21e-06 M=1
+ sca=0.830452 scb=0.000155147 scc=2.70413e-07 lpccnr=2.29e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.215e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XX286/X73/X8/D0_noxref VSS VDD diodenwx  AREA=4.11324e-11 perim=2.72e-05
+ sizedup=0
XXI1/XI5/XI0A/M5P XI1/XI5/XI0A/N3N XI1/XI5/XI0A/N2P VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=7.53851
+ scb=0.00589959 scc=0.000336008 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.05e-07 sb=9.15e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M5P@2 XI1/XI5/XI0A/N3N XI1/XI5/XI0A/N2P VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=7.27107
+ scb=0.00581659 scc=0.00033599 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=3.75e-07 sb=6.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M4P XI1/XI5/XI0A/N2P XI1/XI5/XI0A/N2P VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.24568
+ scb=0.0057654 scc=0.000335987 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=6.45e-07 sb=3.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M4P@2 XI1/XI5/XI0A/N2P XI1/XI5/XI0A/N2P VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=6.24568
+ scb=0.0057654 scc=0.000335987 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=9.15e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M14P XI1/XI5/XI0A/N1N422 XI1/XI5/XI0A/N1N422 VDD VDD pfet
+ L=1.8e-07 W=2e-06 AD=1.2e-13 AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1
+ sca=3.38053 scb=0.00159701 scc=1.61519e-05 lpccnr=1.66e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.05e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M14P@2 XI1/XI5/XI0A/N1N422 XI1/XI5/XI0A/N1N422 VDD VDD pfet
+ L=1.8e-07 W=2e-06 AD=1.2e-13 AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1
+ sca=3.38053 scb=0.00159701 scc=1.61519e-05 lpccnr=1.66e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M14N XI1/XI5/O1 XI1/XI5/XI0A/N1N422 VDD VDD pfet L=1.8e-07 W=2e-06
+ AD=1.2e-13 AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1 sca=3.38053 scb=0.00159701
+ scc=1.61519e-05 lpccnr=1.66e-07 covpccnr=0 wrxcnr=1.8e-06 sa=1.05e-07
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M14N@2 XI1/XI5/O1 XI1/XI5/XI0A/N1N422 VDD VDD pfet L=1.8e-07
+ W=2e-06 AD=1.2e-13 AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1 sca=3.38053
+ scb=0.00159701 scc=1.61519e-05 lpccnr=1.66e-07 covpccnr=0 wrxcnr=1.8e-06
+ sa=4.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M4N XI1/XI5/XI0A/N2N XI1/XI5/XI0A/N2N VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=6.24568
+ scb=0.0057654 scc=0.000335987 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=1.05e-07 sb=9.15e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M4N@2 XI1/XI5/XI0A/N2N XI1/XI5/XI0A/N2N VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=6.24568
+ scb=0.0057654 scc=0.000335987 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=3.75e-07 sb=6.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M5N XI1/XI5/XI0A/N3P XI1/XI5/XI0A/N2N VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=2.124e-13 PD=3.66e-06 PS=3.66e-06 M=1 sca=7.27107
+ scb=0.00581659 scc=0.00033599 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=6.45e-07 sb=3.75e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M5N@2 XI1/XI5/XI0A/N3P XI1/XI5/XI0A/N2N VDD VDD pfet L=1.5e-07
+ W=3.54e-06 AD=2.124e-13 AS=3.717e-13 PD=3.66e-06 PS=7.29e-06 M=1 sca=7.53851
+ scb=0.00589959 scc=0.000336008 lpccnr=1.39e-07 covpccnr=0 wrxcnr=3.186e-06
+ sa=9.15e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0B/MDC3 VDDHA_RX IBRX2 VDDHA_RX VDDHA_RX egpfet L=2e-06 W=6e-06
+ AD=7.2e-13 AS=7.2e-13 PD=1.224e-05 PS=1.224e-05 M=1 sca=4 scb=0.00306566
+ scc=0.000422923 lpccnr=1.815e-06 covpccnr=0 wrxcnr=5.4e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/X1I291/M1 XI1/XI5/XI0A/PDB XI1/PDI VDDHA_RX VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=1.70503 scb=0.000376785 scc=2.23221e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M11P XI1/XI5/XI0A/N2P XI1/XI5/XI0A/PDB VDD VDD egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=18.5703
+ scb=0.0243185 scc=0.000992376 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M1I437 XI1/XI5/XI0A/N1N422 XI1/XI5/XI0A/PDB VDD VDD egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=16.5926 scb=0.0212421 scc=0.000750386 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M1P XI1/XI5/XI0A/N1N IBRX2 XI1/XI5/XI0A/N0 VDDHA_RX egpfet L=3e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0@12 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=5.4e-07 sb=1.8e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0@11 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=9.6e-07 sb=1.38e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M1P@4 XI1/XI5/XI0A/N1N IBRX2 XI1/XI5/XI0A/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=5.6e-07 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0@10 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.38e-06 sb=9.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M1P@3 XI1/XI5/XI0A/N1N IBRX2 XI1/XI5/XI0A/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0@9 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.8e-06 sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M1P@2 XI1/XI5/XI0A/N1N IBRX2 XI1/XI5/XI0A/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.44e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0@8 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0@7 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M1N XI1/XI5/XI0A/N1P XI1/INPI XI1/XI5/XI0A/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0@6 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=5.4e-07 sb=1.8e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M1N@4 XI1/XI5/XI0A/N1P XI1/INPI XI1/XI5/XI0A/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=5.6e-07 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0@5 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=9.6e-07 sb=1.38e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0@4 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.38e-06 sb=9.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M1N@3 XI1/XI5/XI0A/N1P XI1/INPI XI1/XI5/XI0A/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0@3 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.12e-13 PD=1.74e-06 PS=1.74e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.8e-06 sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M1N@2 XI1/XI5/XI0A/N1P XI1/INPI XI1/XI5/XI0A/N0 VDDHA_RX egpfet
+ L=3e-07 W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.44e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M0@2 XI1/XI5/XI0A/N0 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=4.40381
+ scb=0.00434195 scc=0.000147722 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M11N XI1/XI5/XI0A/N2N XI1/XI5/XI0A/PDB VDD VDD egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=18.5703
+ scb=0.0243185 scc=0.000992376 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M7N XI1/XI5/XI0A/N3N XI1/XI5/XI0A/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=1.005e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0A/M7N@2 XI1/XI5/XI0A/N3N XI1/XI5/XI0A/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=4.05e-07 sb=7.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0A/M6P XI1/XI5/XI0A/N3N XI1/XI5/XI0A/N3N VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=7.05e-07 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0A/M6P@2 XI1/XI5/XI0A/N3N XI1/XI5/XI0A/N3N VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.005e-06 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0A/M13P XI1/XI5/XI0A/N1N422 XI1/XI5/XI0A/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0A/M13P@2 XI1/XI5/XI0A/N1N422 XI1/XI5/XI0A/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=4.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0A/M10P XI1/XI5/XI0A/N3N XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M12P XI1/XI5/XI0A/N1N XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M7P XI1/XI5/XI0A/N3P XI1/XI5/XI0A/N3N VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=1.005e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0A/M7P@2 XI1/XI5/XI0A/N3P XI1/XI5/XI0A/N3N VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=4.05e-07 sb=7.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0A/M6N XI1/XI5/XI0A/N3P XI1/XI5/XI0A/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=7.05e-07 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0A/M6N@2 XI1/XI5/XI0A/N3P XI1/XI5/XI0A/N3P VSSA_RX VSSA_RX nfet
+ L=1.8e-07 W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.005e-06 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0A/M13N XI1/XI5/O1 XI1/XI5/XI0A/N3N VSSA_RX VSSA_RX nfet L=1.8e-07
+ W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=4.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M13N@2 XI1/XI5/O1 XI1/XI5/XI0A/N3N VSSA_RX VSSA_RX nfet L=1.8e-07
+ W=1e-06 AD=6e-14 AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.66e-07 covpccnr=0 wrxcnr=9e-07 sa=4.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M10N XI1/XI5/XI0A/N3P XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/M12N XI1/XI5/XI0A/N1P XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XI0A/X1I291/M2 XI1/XI5/XI0A/PDB XI1/PDI VSSA_RX VSSA_RX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XI0A/M13 XI1/XI5/O1 XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC0@22 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=6e-13
+ PD=5.14e-06 PS=1.024e-05 M=1 sca=2.17718 scb=0.00103367 scc=1.0163e-05
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@21 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@20 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@19 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@18 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@17 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@16 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=6e-13 AS=3.5e-13
+ PD=1.024e-05 PS=5.14e-06 M=1 sca=2.17718 scb=0.00103367 scc=1.0163e-05
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI3/X1I124/M0 XI1/XI3/TIEL XI1/XI3/X1I124/N1N50 VSS VSS nfet L=3e-08
+ W=1.1e-07 AD=2.09e-14 AS=2.09e-14 PD=6e-07 PS=6e-07 M=1 sca=3.38327
+ scb=0.000920314 scc=1.06271e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9.9e-08
+ sa=1.9e-07 sb=1.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC0@15 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=6e-13
+ PD=5.14e-06 PS=1.024e-05 M=1 sca=2.17718 scb=0.00103367 scc=1.0163e-05
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@14 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@13 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@12 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@11 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@10 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@9 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=6e-13 AS=3.5e-13
+ PD=1.024e-05 PS=5.14e-06 M=1 sca=2.17718 scb=0.00103367 scc=1.0163e-05
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI3/X1I124/M1 XI1/XI3/X1I124/N1N50 XI1/XI3/X1I124/N1N50 VDD VDD pfet
+ L=3e-08 W=1.1e-07 AD=2.09e-14 AS=2.09e-14 PD=6e-07 PS=6e-07 M=1 sca=109.038
+ scb=0.0600072 scc=0.0149457 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9.9e-08
+ sa=1.9e-07 sb=1.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC0@8 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=6e-13
+ PD=5.14e-06 PS=1.024e-05 M=1 sca=2.17718 scb=0.00103367 scc=1.0163e-05
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@7 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@6 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@5 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@4 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@3 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=3.5e-13 AS=3.5e-13
+ PD=5.14e-06 PS=5.14e-06 M=1 sca=1.14755 scb=0.000590218 scc=6.64827e-06
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC0@2 VDD VSS VDD VDD egpfet L=5e-06 W=5e-06 AD=6e-13 AS=3.5e-13
+ PD=1.024e-05 PS=5.14e-06 M=1 sca=2.17718 scb=0.00103367 scc=1.0163e-05
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC2@15 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@14 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@13 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@12 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG7A/M2 XI1/XI3/N4A XI1/XI3/N3A VSS VSS nfet L=3e-08 W=1.26e-06
+ AD=1.323e-13 AS=1.323e-13 PD=2.73e-06 PS=2.73e-06 M=1 sca=0.771574
+ scb=2.1376e-05 scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG8A/M2 XI1/XI3/N5A XI1/XI3/N4A VSS VSS nfet L=3e-08 W=1.26e-06
+ AD=7.56e-14 AS=1.323e-13 PD=1.38e-06 PS=2.73e-06 M=1 sca=0.771574
+ scb=2.1376e-05 scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06
+ sa=1.05e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG8A/M2@3 XI1/XI3/N5A XI1/XI3/N4A VSS VSS nfet L=3e-08 W=1.26e-06
+ AD=7.56e-14 AS=7.56e-14 PD=1.38e-06 PS=1.38e-06 M=1 sca=0.771574
+ scb=2.1376e-05 scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06
+ sa=2.55e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG8A/M2@2 XI1/XI3/N5A XI1/XI3/N4A VSS VSS nfet L=3e-08 W=1.26e-06
+ AD=1.323e-13 AS=7.56e-14 PD=2.73e-06 PS=1.38e-06 M=1 sca=0.771574
+ scb=2.1376e-05 scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06
+ sa=4.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M2 DOI XI1/XI3/N5A VSS VSS nfet L=3e-08 W=1.26e-06 AD=7.56e-14
+ AS=1.323e-13 PD=1.38e-06 PS=2.73e-06 M=1 sca=0.771574 scb=2.1376e-05
+ scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06 sa=1.05e-07
+ sb=1.305e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M2@9 DOI XI1/XI3/N5A VSS VSS nfet L=3e-08 W=1.26e-06 AD=7.56e-14
+ AS=7.56e-14 PD=1.38e-06 PS=1.38e-06 M=1 sca=0.771574 scb=2.1376e-05
+ scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06 sa=2.55e-07
+ sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M2@8 DOI XI1/XI3/N5A VSS VSS nfet L=3e-08 W=1.26e-06 AD=7.56e-14
+ AS=7.56e-14 PD=1.38e-06 PS=1.38e-06 M=1 sca=0.771574 scb=2.1376e-05
+ scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06 sa=4.05e-07
+ sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M2@7 DOI XI1/XI3/N5A VSS VSS nfet L=3e-08 W=1.26e-06 AD=7.56e-14
+ AS=7.56e-14 PD=1.38e-06 PS=1.38e-06 M=1 sca=0.771574 scb=2.1376e-05
+ scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06 sa=5.55e-07
+ sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M2@6 DOI XI1/XI3/N5A VSS VSS nfet L=3e-08 W=1.26e-06 AD=7.56e-14
+ AS=7.56e-14 PD=1.38e-06 PS=1.38e-06 M=1 sca=0.771574 scb=2.1376e-05
+ scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06 sa=7.05e-07
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M2@5 DOI XI1/XI3/N5A VSS VSS nfet L=3e-08 W=1.26e-06 AD=7.56e-14
+ AS=7.56e-14 PD=1.38e-06 PS=1.38e-06 M=1 sca=0.771574 scb=2.1376e-05
+ scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06 sa=8.55e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M2@4 DOI XI1/XI3/N5A VSS VSS nfet L=3e-08 W=1.26e-06 AD=7.56e-14
+ AS=7.56e-14 PD=1.38e-06 PS=1.38e-06 M=1 sca=0.771574 scb=2.1376e-05
+ scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06 sa=1.005e-06
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M2@3 DOI XI1/XI3/N5A VSS VSS nfet L=3e-08 W=1.26e-06 AD=7.56e-14
+ AS=7.56e-14 PD=1.38e-06 PS=1.38e-06 M=1 sca=0.771574 scb=2.1376e-05
+ scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06 sa=1.155e-06
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M2@2 DOI XI1/XI3/N5A VSS VSS nfet L=3e-08 W=1.26e-06 AD=1.323e-13
+ AS=7.56e-14 PD=2.73e-06 PS=1.38e-06 M=1 sca=0.771574 scb=2.1376e-05
+ scc=1.10074e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.134e-06 sa=1.305e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG7A/M1 XI1/XI3/N4A XI1/XI3/N3A VDD VDD pfet L=3e-08 W=2.9e-06
+ AD=3.045e-13 AS=3.045e-13 PD=6.01e-06 PS=6.01e-06 M=1 sca=10.4885
+ scb=0.00708963 scc=0.0010505 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.61e-06
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG8A/M1 XI1/XI3/N5A XI1/XI3/N4A VDD VDD pfet L=3e-08 W=2.52e-06
+ AD=1.512e-13 AS=2.646e-13 PD=2.64e-06 PS=5.25e-06 M=1 sca=11.522
+ scb=0.00790192 scc=0.00120804 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06
+ sa=1.05e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG8A/M1@3 XI1/XI3/N5A XI1/XI3/N4A VDD VDD pfet L=3e-08 W=2.52e-06
+ AD=1.512e-13 AS=1.512e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=11.522
+ scb=0.00790192 scc=0.00120804 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06
+ sa=2.55e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI3/XG8A/M1@2 XI1/XI3/N5A XI1/XI3/N4A VDD VDD pfet L=3e-08 W=2.52e-06
+ AD=2.646e-13 AS=1.512e-13 PD=5.25e-06 PS=2.64e-06 M=1 sca=12.5301 scb=0.007949
+ scc=0.00120804 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06 sa=4.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M1 DOI XI1/XI3/N5A VDD VDD pfet L=3e-08 W=2.52e-06 AD=1.512e-13
+ AS=2.646e-13 PD=2.64e-06 PS=5.25e-06 M=1 sca=13.4728 scb=0.00845853
+ scc=0.00120848 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06 sa=1.05e-07
+ sb=1.305e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M1@9 DOI XI1/XI3/N5A VDD VDD pfet L=3e-08 W=2.52e-06 AD=1.512e-13
+ AS=1.512e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=13.846 scb=0.00883112
+ scc=0.00120936 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06 sa=2.55e-07
+ sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M1@8 DOI XI1/XI3/N5A VDD VDD pfet L=3e-08 W=2.52e-06 AD=1.512e-13
+ AS=1.512e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=14.3375 scb=0.00944016
+ scc=0.00121202 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06 sa=4.05e-07
+ sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M1@7 DOI XI1/XI3/N5A VDD VDD pfet L=3e-08 W=2.52e-06 AD=1.512e-13
+ AS=1.512e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=15.0032 scb=0.0104225
+ scc=0.00121991 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06 sa=5.55e-07
+ sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M1@6 DOI XI1/XI3/N5A VDD VDD pfet L=3e-08 W=2.52e-06 AD=1.512e-13
+ AS=1.512e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=15.9362 scb=0.0119806
+ scc=0.00124303 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06 sa=7.05e-07
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M1@5 DOI XI1/XI3/N5A VDD VDD pfet L=3e-08 W=2.52e-06 AD=1.512e-13
+ AS=1.512e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=17.3017 scb=0.0143967
+ scc=0.00130956 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06 sa=8.55e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M1@4 DOI XI1/XI3/N5A VDD VDD pfet L=3e-08 W=2.52e-06 AD=1.512e-13
+ AS=1.512e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=19.4147 scb=0.0180288
+ scc=0.00149646 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06 sa=1.005e-06
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M1@3 DOI XI1/XI3/N5A VDD VDD pfet L=3e-08 W=2.52e-06 AD=1.512e-13
+ AS=1.512e-13 PD=2.64e-06 PS=2.64e-06 M=1 sca=22.9401 scb=0.0232433
+ scc=0.00200412 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06 sa=1.155e-06
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI3/XG9A/M1@2 DOI XI1/XI3/N5A VDD VDD pfet L=3e-08 W=2.52e-06 AD=2.646e-13
+ AS=1.512e-13 PD=5.25e-06 PS=2.64e-06 M=1 sca=29.4882 scb=0.0301871
+ scc=0.00331493 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.268e-06 sa=1.305e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XX286/X88/D0_noxref VSS VDD diodenwx  AREA=1.66314e-11 perim=1.663e-05 sizedup=0
XXI1/XI5/RR0 VSSA_RX XI1/XI5/N1N312 VDDHA_RX opppcres 1701.34 M=1 w=2e-06
+ l=5.51e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/XG2/M2 XI1/VAL XI1/XI5/N1N356 VSS VSS nfet L=3e-08 W=1.8e-06
+ AD=1.89e-13 AS=1.89e-13 PD=3.81e-06 PS=3.81e-06 M=1 sca=1.00176
+ scb=9.94212e-05 scc=4.17215e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XG1/M2 XI1/XI5/N1N356 XI1/XI5/N1N284 VSS VSS nfet L=3e-08 W=9e-07
+ AD=9.45e-14 AS=9.45e-14 PD=2.01e-06 PS=2.01e-06 M=1 sca=1.34134
+ scb=0.000191241 scc=8.33511e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=8.1e-07
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XG0/M4 XI1/XI5/XG0/N1 XI1/XI5/O2 VSS VSS nfet L=3e-08 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=1.29265 scb=0.000174293
+ scc=7.50603e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=2.55e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XG0/M3 XI1/XI5/N1N284 XI1/XI5/O1 XI1/XI5/XG0/N1 VSS nfet L=3e-08
+ W=1e-06 AD=1.05e-13 AS=6e-14 PD=2.21e-06 PS=1.12e-06 M=1 sca=1.29265
+ scb=0.000174293 scc=7.50603e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07
+ sa=2.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI5/XG2/M1 XI1/VAL XI1/XI5/N1N356 VDD VDD pfet L=3e-08 W=3.6e-06
+ AD=3.78e-13 AS=3.78e-13 PD=7.41e-06 PS=7.41e-06 M=1 sca=14.331 scb=0.0168296
+ scc=0.000672162 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI5/XG1/M1 XI1/XI5/N1N356 XI1/XI5/N1N284 VDD VDD pfet L=3e-08 W=1.8e-06
+ AD=1.89e-13 AS=1.89e-13 PD=3.81e-06 PS=3.81e-06 M=1 sca=10.2544 scb=0.00820741
+ scc=0.000126429 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI5/XG0/M2 XI1/XI5/N1N284 XI1/XI5/O2 VDD VDD pfet L=3e-08 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=10.4314 scb=0.00881986
+ scc=0.000144303 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=2.55e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/XG0/M1 XI1/XI5/N1N284 XI1/XI5/O1 VDD VDD pfet L=3e-08 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=11.5164 scb=0.0109676
+ scc=0.000198226 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=2.55e-07 sb=1.05e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI5/RRD3 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 8306.07 M=1 w=1e-06
+ l=1.356e-05   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/RRD4 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 8306.07 M=1 w=1e-06
+ l=1.356e-05   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/RR5 IBRX2 IBRX2 VDDHA_RX opppcres 467.791 M=1 w=1.46e-06 l=1e-06   bp=1
+ pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/RR6 IBRX2 IBRX2 VDDHA_RX opppcres 467.791 M=1 w=1.46e-06 l=1e-06   bp=1
+ pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/RR7 IBRX2 IBRX2 VDDHA_RX opppcres 467.791 M=1 w=1.46e-06 l=1e-06   bp=1
+ pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/RR8 IBRX2 IBRX2 VDDHA_RX opppcres 467.791 M=1 w=1.46e-06 l=1e-06   bp=1
+ pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/RR1 XI1/XI5/N1N312 X286/X88/noxref_55 VDDHA_RX opppcres 467.791 M=1
+ w=1.46e-06 l=1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/RR2 X286/X88/noxref_55 X286/X88/noxref_56 VDDHA_RX opppcres 467.791 M=1
+ w=1.46e-06 l=1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/RR3 X286/X88/noxref_56 X286/X88/noxref_57 VDDHA_RX opppcres 467.791 M=1
+ w=1.46e-06 l=1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/RR4 X286/X88/noxref_57 IBRX2 VDDHA_RX opppcres 467.791 M=1 w=1.46e-06
+ l=1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/RRD1 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 4641.35 M=1 w=1e-06 l=7.52e-06
+ bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI1/XI5/RRD2 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 4641.35 M=1 w=1e-06 l=7.52e-06
+ bp=1 pbar=1 s=1 ncr=1 sizedup=0
XX286/X89/D0_noxref VSS VDD diodenwx  AREA=5.39748e-11 perim=3.122e-05 sizedup=0
XXI1/XI4/M6N XI1/NN XI1/INP2 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14 AS=1.05e-13
+ PD=1.12e-06 PS=2.21e-06 M=1 sca=0.912112 scb=4.07878e-05 scc=3.44045e-09
+ lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=1.645e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M6N@2 XI1/NN XI1/INP2 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14 AS=6e-14
+ PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05 scc=3.44045e-09
+ lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=3.25e-07 sb=1.425e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M5N XI1/NN XI1/INP1 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14 AS=6e-14
+ PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05 scc=3.44045e-09
+ lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=5.45e-07 sb=1.205e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M5N@2 XI1/NN XI1/INP1 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14 AS=6e-14
+ PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05 scc=3.44045e-09
+ lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=7.65e-07 sb=9.85e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M6P XI1/XI4/N1N XI1/INN2 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14 AS=6e-14
+ PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05 scc=3.44045e-09
+ lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=9.85e-07 sb=7.65e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M6P@2 XI1/XI4/N1N XI1/INN2 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05
+ scc=3.44045e-09 lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=1.205e-06
+ sb=5.45e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M5P XI1/XI4/N1N XI1/INN1 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14 AS=6e-14
+ PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05 scc=3.44045e-09
+ lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=1.425e-06 sb=3.25e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M5P@2 XI1/XI4/N1N XI1/INN1 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0.912112 scb=4.07878e-05
+ scc=3.44045e-09 lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=1.645e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M1P XI1/XI4/N1P XI1/INP1 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0.912112 scb=4.07878e-05
+ scc=3.44045e-09 lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07
+ sb=1.645e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M1P@2 XI1/XI4/N1P XI1/INP1 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05
+ scc=3.44045e-09 lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=3.25e-07
+ sb=1.425e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M2P XI1/XI4/N1P XI1/INP2 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14 AS=6e-14
+ PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05 scc=3.44045e-09
+ lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=5.45e-07 sb=1.205e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M2P@2 XI1/XI4/N1P XI1/INP2 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05
+ scc=3.44045e-09 lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=7.65e-07 sb=9.85e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI4/M1N XI1/NP XI1/INN1 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14 AS=6e-14
+ PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05 scc=3.44045e-09
+ lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=9.85e-07 sb=7.65e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M1N@2 XI1/NP XI1/INN1 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14 AS=6e-14
+ PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05 scc=3.44045e-09
+ lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=1.205e-06 sb=5.45e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M2N XI1/NP XI1/INN2 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14 AS=6e-14
+ PD=1.12e-06 PS=1.12e-06 M=1 sca=0.912112 scb=4.07878e-05 scc=3.44045e-09
+ lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=1.425e-06 sb=3.25e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M2N@2 XI1/NP XI1/INN2 VSS VSS nfet L=1e-07 W=1e-06 AD=6e-14 AS=1.05e-13
+ PD=1.12e-06 PS=2.21e-06 M=1 sca=0.912112 scb=4.07878e-05 scc=3.44045e-09
+ lpccnr=9.4e-08 covpccnr=0 wrxcnr=9e-07 sa=1.645e-06 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M1 XI1/NP XI1/PDI VSS VSS egnfet L=1.5e-07 W=4e-07 AD=4.8e-14
+ AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=1.68726 scb=0.000363943
+ scc=2.07183e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI4/X1I229/M2 XI1/XI4/PDB XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI4/M4N XI1/NN XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1 sca=4.63009 scb=0.00245123
+ scc=4.89204e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.05e-07
+ sb=2.0022e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M4N@6 XI1/NN XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=3.05e-07
+ sb=2.0022e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M4N@5 XI1/NN XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=5.05e-07
+ sb=1.905e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M4N@4 XI1/NN XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=7.05e-07
+ sb=1.705e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M4N@3 XI1/NN XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=9.05e-07
+ sb=1.505e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M4N@2 XI1/NN XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.105e-06
+ sb=1.305e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M4P XI1/XI4/N1N XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.305e-06
+ sb=1.105e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M4P@6 XI1/XI4/N1N XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.505e-06
+ sb=9.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M4P@5 XI1/XI4/N1N XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.705e-06
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M4P@4 XI1/XI4/N1N XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.905e-06
+ sb=5.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M4P@3 XI1/XI4/N1N XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=2.0022e-06
+ sb=3.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M4P@2 XI1/XI4/N1N XI1/XI4/N1N VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=2.0022e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3P XI1/XI4/N1P XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.05e-07
+ sb=2.0022e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3P@6 XI1/XI4/N1P XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=3.05e-07
+ sb=2.0022e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3P@5 XI1/XI4/N1P XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=5.05e-07
+ sb=1.905e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3P@4 XI1/XI4/N1P XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=7.05e-07
+ sb=1.705e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3P@3 XI1/XI4/N1P XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=9.05e-07
+ sb=1.505e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3P@2 XI1/XI4/N1P XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.105e-06
+ sb=1.305e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3N XI1/NP XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.305e-06
+ sb=1.105e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3N@6 XI1/NP XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.505e-06
+ sb=9.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3N@5 XI1/NP XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.705e-06
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3N@4 XI1/NP XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.905e-06
+ sb=5.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3N@3 XI1/NP XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=1.2e-13 PD=2.12e-06 PS=2.12e-06 M=1 sca=3.54472 scb=0.00238599
+ scc=4.89159e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=2.0022e-06
+ sb=3.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M3N@2 XI1/NP XI1/XI4/N1P VDD VDD pfet L=8e-08 W=2e-06 AD=1.2e-13
+ AS=2.1e-13 PD=2.12e-06 PS=4.21e-06 M=1 sca=4.63009 scb=0.00245123
+ scc=4.89204e-05 lpccnr=7.6e-08 covpccnr=0 wrxcnr=1.8e-06 sa=2.0022e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI4/M2 XI1/NN XI1/XI4/PDB VDD VDD egpfet L=1.5e-07 W=4e-07 AD=4.8e-14
+ AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=15.6288 scb=0.0198062
+ scc=0.000611806 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI4/M1I308 XI1/XI4/N1N XI1/XI4/PDB VDD VDD egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=9.88869 scb=0.0113889
+ scc=0.000381701 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI4/M1I225 XI1/XI4/N1P XI1/XI4/PDB VDD VDD egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=12.25 scb=0.0140798
+ scc=0.000302066 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI4/X1I229/M1 XI1/XI4/PDB XI1/PDI VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=4.62809
+ scb=0.00269551 scc=1.33705e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/M4N XI1/XI6/N3 PDRXI VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=3.07821 scb=0.00190794
+ scc=6.39406e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI6/XG2/M2 XI1/PDI XI1/XI6/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/XG2/M2@4 XI1/PDI XI1/XI6/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/XG2/M2@3 XI1/PDI XI1/XI6/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/XG2/M2@2 XI1/PDI XI1/XI6/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/XG1/M2 XI1/XI6/N1N36 XI1/XI6/N1N5 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/M4P XI1/XI6/N1N5 XI1/XI6/N2 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/M3N XI1/XI6/N3 PDRXI VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=29.0407 scb=0.033526
+ scc=0.00176982 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI6/XG2/M1 XI1/PDI XI1/XI6/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=9.42555
+ scb=0.0100427 scc=0.000276867 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/XG2/M1@4 XI1/PDI XI1/XI6/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=7.10155
+ scb=0.00601223 scc=0.000177513 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/XG2/M1@3 XI1/PDI XI1/XI6/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=5.91934
+ scb=0.00433708 scc=0.000164871 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/XG2/M1@2 XI1/PDI XI1/XI6/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=5.23693
+ scb=0.00368289 scc=0.000163346 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/XG1/M1 XI1/XI6/N1N36 XI1/XI6/N1N5 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=3.36e-13 AS=3.36e-13 PD=5.84e-06 PS=5.84e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/M3P XI1/XI6/N1N5 XI1/XI6/N2 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=3.43331
+ scb=0.00285132 scc=4.77845e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/M1P XI1/XI6/N2 XI1/XI6/N1 VDDHA_RX VDDHA_RX egpfet L=3e-06 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979 scb=0.00151603
+ scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI6/M1N XI1/XI6/N1 XI1/XI6/N2 VDDHA_RX VDDHA_RX egpfet L=3e-06 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=4.11762 scb=0.0021369
+ scc=3.00661e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI6/M2P XI1/XI6/N2 PDRXI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI6/M2N XI1/XI6/N1 XI1/XI6/N3 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1N XI1/XI2/N1N XI1/INPI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1N@6 XI1/XI2/N1N XI1/INPI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=6.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1N@5 XI1/XI2/N1N XI1/INPI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.1e-06 sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1N@4 XI1/XI2/N1N XI1/INPI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.59e-06 sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1N@3 XI1/XI2/N1N XI1/INPI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=2.0083e-06 sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1N@2 XI1/XI2/N1N XI1/INPI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1P XI1/XI2/N1P XI1/INNI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1P@6 XI1/XI2/N1P XI1/INNI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=6.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1P@5 XI1/XI2/N1P XI1/INNI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.1e-06 sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1P@4 XI1/XI2/N1P XI1/INNI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.59e-06 sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1P@3 XI1/XI2/N1P XI1/INNI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=2.0083e-06 sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M1P@2 XI1/XI2/N1P XI1/INNI XI1/XI2/N1N204 VSSA_RX egnfet L=3.5e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0.464215
+ scb=1.86788e-05 scc=3.75552e-09 lpccnr=3.3e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/X1I277/M1 XI1/XI2/PDIB XI1/PDI VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=9.15751
+ scb=0.011838 scc=0.00050139 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/X1I279/M1 XI1/XI2/PDI XI1/XI2/PDIB VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=9.15751
+ scb=0.011838 scc=0.00050139 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/X1I277/M2 XI1/XI2/PDIB XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/X1I279/M2 XI1/XI2/PDI XI1/XI2/PDIB VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M4N XI1/INP2 XI1/INP2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=1.645e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M4N@4 XI1/INP2 XI1/INP2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=3.25e-07 sb=1.425e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M4N@3 XI1/INP2 XI1/INP2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=5.45e-07 sb=1.205e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M4N@2 XI1/INP2 XI1/INP2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=7.65e-07 sb=9.85e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M5P XI1/INP2 XI1/INN2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=9.85e-07 sb=7.65e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M5P@4 XI1/INP2 XI1/INN2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.205e-06 sb=5.45e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M5P@3 XI1/INP2 XI1/INN2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.425e-06 sb=3.25e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M5P@2 XI1/INP2 XI1/INN2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.645e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M0 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=1.44e-13 PD=1.34e-06 PS=2.64e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@24 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=5.6e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M9N XI1/INP2 XI1/XI2/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M0@23 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@22 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.44e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@21 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.88e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@20 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@19 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@18 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=1.88e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@17 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=1.44e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@16 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=1e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@15 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=5.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@14 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=1.44e-13 PD=1.34e-06 PS=2.64e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M2N XI1/XI2/N1N XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI2/M2N@6 XI1/XI2/N1N XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.5e-06 AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436
+ scb=9.4701e-05 scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06
+ sa=5.6e-07 sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M2N@5 XI1/XI2/N1N XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.5e-06 AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436
+ scb=9.4701e-05 scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06
+ sa=1e-06 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M2N@4 XI1/XI2/N1N XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.5e-06 AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436
+ scb=9.4701e-05 scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06
+ sa=1.44e-06 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M2N@3 XI1/XI2/N1N XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.5e-06 AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436
+ scb=9.4701e-05 scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06
+ sa=1.88e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M2N@2 XI1/XI2/N1N XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1 sca=1.03436
+ scb=9.4701e-05 scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M3N XI1/INP2 XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI2/M3N@6 XI1/INP2 XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=5.6e-07
+ sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI2/M3N@5 XI1/INP2 XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=1e-06 sb=1.44e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M3N@4 XI1/INP2 XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=1.44e-06 sb=1e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M3N@3 XI1/INP2 XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=1.88e-06
+ sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI2/M3N@2 XI1/INP2 XI1/XI2/N1N VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI2/M8N XI1/XI2/N1N XI1/XI2/PDIB VDDHA_RX VDDHA_RX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M4P XI1/INN2 XI1/INN2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=1.645e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M4P@4 XI1/INN2 XI1/INN2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=3.25e-07 sb=1.425e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M4P@3 XI1/INN2 XI1/INN2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=5.45e-07 sb=1.205e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M4P@2 XI1/INN2 XI1/INN2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=7.65e-07 sb=9.85e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M5N XI1/INN2 XI1/INP2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=9.85e-07 sb=7.65e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M5N@4 XI1/INN2 XI1/INP2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.205e-06 sb=5.45e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M5N@3 XI1/INN2 XI1/INP2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=6e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.425e-06 sb=3.25e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M5N@2 XI1/INN2 XI1/INP2 VSSA_RX VSSA_RX nfet L=1e-07 W=1e-06 AD=6e-14
+ AS=1.05e-13 PD=1.12e-06 PS=2.21e-06 M=1 sca=0 scb=0 scc=0 lpccnr=9.4e-08
+ covpccnr=0 wrxcnr=9e-07 sa=1.645e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M0@13 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=1.44e-13 PD=1.34e-06 PS=2.64e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@12 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=5.6e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M9P XI1/INN2 XI1/XI2/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M0@11 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@10 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.44e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@9 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.88e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@8 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@7 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@6 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=1.88e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@5 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=1.44e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@4 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=1e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@3 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=8.4e-14 PD=1.34e-06 PS=1.34e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=5.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M0@2 XI1/XI2/N1N204 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=1.44e-13 PD=1.34e-06 PS=2.64e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M2P XI1/XI2/N1P XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI2/M2P@6 XI1/XI2/N1P XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.5e-06 AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436
+ scb=9.4701e-05 scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06
+ sa=5.6e-07 sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M2P@5 XI1/XI2/N1P XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.5e-06 AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436
+ scb=9.4701e-05 scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06
+ sa=1e-06 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M2P@4 XI1/XI2/N1P XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.5e-06 AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436
+ scb=9.4701e-05 scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06
+ sa=1.44e-06 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M2P@3 XI1/XI2/N1P XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.5e-06 AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436
+ scb=9.4701e-05 scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06
+ sa=1.88e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M2P@2 XI1/XI2/N1P XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1 sca=1.03436
+ scb=9.4701e-05 scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI2/M3P XI1/INN2 XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI2/M3P@6 XI1/INN2 XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=5.6e-07
+ sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI2/M3P@5 XI1/INN2 XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=1e-06 sb=1.44e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M3P@4 XI1/INN2 XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=1.44e-06 sb=1e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI2/M3P@3 XI1/INN2 XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=1.88e-06
+ sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI2/M3P@2 XI1/INN2 XI1/XI2/N1P VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.5e-06
+ AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1 sca=1.03436 scb=9.4701e-05
+ scc=3.0794e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.35e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI2/M8P XI1/XI2/N1P XI1/XI2/PDIB VDDHA_RX VDDHA_RX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/MDC1 VSSA_RX XI1/XI0/N7 VSSA_RX VSSA_RX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI0/MDC1@2 VSSA_RX XI1/XI0/N7 VSSA_RX VSSA_RX egnfet L=5e-06 W=5e-06
+ AD=6e-13 AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI0/X1I117/M2 XI1/XI0/PDB XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M15 XI1/XI0/N8 XI1/XI0/N7 VSSA_RX VSSA_RX egnfet L=6e-07 W=7.4e-07
+ AD=8.88e-14 AS=8.88e-14 PD=1.72e-06 PS=1.72e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=5.55e-07 covpccnr=0 wrxcnr=6.66e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M18 XI1/VBN XI1/XI0/N7 XI1/XI0/N10 VSSA_RX egnfet L=3e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07 sb=5.6e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M18@2 XI1/VBN XI1/XI0/N7 XI1/XI0/N10 VSSA_RX egnfet L=3e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=2.16e-06 sa=5.6e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/MDC3 VDDHA_RX XI1/XI0/N2 VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=12.9662 scb=0.0103862
+ scc=0.00132133 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI0/MDC3@2 VDDHA_RX XI1/XI0/N2 VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=9.52381 scb=0.00735759
+ scc=0.00101501 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI0/X1I117/M1 XI1/XI0/PDB XI1/PDI VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=17.6137
+ scb=0.0228038 scc=0.000868969 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M1I54 XI1/XI0/N2 XI1/XI0/PDB VDDHA_RX VDDHA_RX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=9.39002 scb=0.0121669
+ scc=0.000535984 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI0/M5 XI1/XI0/N2 XI1/XI0/N2 XI1/XI0/N3 VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=0.841683
+ scb=4.07986e-05 scc=5.52866e-09 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=1.2e-07 sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M4 XI1/XI0/N3 XI1/XI0/N2 VDDHA_RX VDDHA_RX egpfet L=3e-07 W=7e-07
+ AD=8.4e-14 AS=8.4e-14 PD=1.64e-06 PS=1.64e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M5@2 XI1/XI0/N2 XI1/XI0/N2 XI1/XI0/N3 VDDHA_RX egpfet L=2.8e-07
+ W=1.6e-06 AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=0.841683
+ scb=4.07986e-05 scc=5.52866e-09 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06
+ sa=5.4e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M9 XI1/VBP XI1/XI0/N2 XI1/XI0/N4 VDDHA_RX egpfet L=2.8e-07 W=3.84e-06
+ AD=2.688e-13 AS=4.608e-13 PD=3.98e-06 PS=7.92e-06 M=1 sca=0.509222
+ scb=1.50469e-05 scc=1.76918e-09 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.456e-06
+ sa=1.2e-07 sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M8 XI1/XI0/N4 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=3.02513 scb=0.00232059
+ scc=3.51389e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=1.2e-07
+ sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI0/M9@2 XI1/VBP XI1/XI0/N2 XI1/XI0/N4 VDDHA_RX egpfet L=2.8e-07 W=3.84e-06
+ AD=2.688e-13 AS=4.608e-13 PD=3.98e-06 PS=7.92e-06 M=1 sca=0.509222
+ scb=1.50469e-05 scc=1.76918e-09 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.456e-06
+ sa=5.4e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M8@2 XI1/XI0/N4 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=3.02513 scb=0.00232059
+ scc=3.51389e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=5.4e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI0/M1I189 XI1/VBP XI1/XI0/PDB VDDHA_RX VDDHA_RX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=9.39002 scb=0.0121669
+ scc=0.000535984 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/XI0/M13 XI1/XI0/N7 XI1/XI0/N2 XI1/XI0/N6 VDDHA_RX egpfet L=2.8e-07
+ W=3.84e-06 AD=2.688e-13 AS=4.608e-13 PD=3.98e-06 PS=7.92e-06 M=1 sca=0.521042
+ scb=1.70475e-05 scc=2.30362e-09 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.456e-06
+ sa=1.2e-07 sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M12 XI1/XI0/N6 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=3.02513 scb=0.00232059
+ scc=3.51389e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=1.2e-07
+ sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI0/M13@2 XI1/XI0/N7 XI1/XI0/N2 XI1/XI0/N6 VDDHA_RX egpfet L=2.8e-07
+ W=3.84e-06 AD=2.688e-13 AS=4.608e-13 PD=3.98e-06 PS=7.92e-06 M=1 sca=0.521042
+ scb=1.70475e-05 scc=2.30362e-09 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.456e-06
+ sa=5.4e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M12@2 XI1/XI0/N6 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=3.02513 scb=0.00232059
+ scc=3.51389e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=5.4e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI0/M16 XI1/XI0/N9 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=3.02513 scb=0.00232059
+ scc=3.51389e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=1.2e-07
+ sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI0/M17 XI1/VBN XI1/XI0/N2 XI1/XI0/N9 VDDHA_RX egpfet L=2.8e-07 W=3.84e-06
+ AD=2.688e-13 AS=4.608e-13 PD=3.98e-06 PS=7.92e-06 M=1 sca=0.521042
+ scb=1.70475e-05 scc=2.30362e-09 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.456e-06
+ sa=1.2e-07 sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M16@2 XI1/XI0/N9 XI1/VBP VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=1.6e-06
+ AD=1.12e-13 AS=1.92e-13 PD=1.74e-06 PS=3.44e-06 M=1 sca=3.02513 scb=0.00232059
+ scc=3.51389e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=1.44e-06 sa=5.4e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/XI0/M17@2 XI1/VBN XI1/XI0/N2 XI1/XI0/N9 VDDHA_RX egpfet L=2.8e-07
+ W=3.84e-06 AD=2.688e-13 AS=4.608e-13 PD=3.98e-06 PS=7.92e-06 M=1 sca=0.521042
+ scb=1.70475e-05 scc=2.30362e-09 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.456e-06
+ sa=5.4e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M1I77 XI1/XI0/N7 XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M1I82 XI1/VBN XI1/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M14 XI1/XI0/N7 XI1/XI0/N7 XI1/XI0/N8 VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=1.44e-13 PD=1.34e-06 PS=2.64e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.2e-07 sb=5.6e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M14@2 XI1/XI0/N7 XI1/XI0/N7 XI1/XI0/N8 VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=1.44e-13 PD=1.34e-06 PS=2.64e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=5.6e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M19 XI1/XI0/N10 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=1.44e-13 PD=1.34e-06 PS=2.64e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.2e-07 sb=5.6e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M19@2 XI1/XI0/N10 XI1/VBN VSSA_RX VSSA_RX egnfet L=3e-07 W=1.2e-06
+ AD=8.4e-14 AS=1.44e-13 PD=1.34e-06 PS=2.64e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.08e-06 sa=5.6e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M3 IBRX1 IBRX1 VSSA_RX VSSA_RX egnfet L=3e-07 W=8e-07 AD=5.6e-14
+ AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M3@2 IBRX1 IBRX1 VSSA_RX VSSA_RX egnfet L=3e-07 W=8e-07 AD=5.6e-14
+ AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=5.6e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M7 XI1/XI0/N2 IBRX1 VSSA_RX VSSA_RX egnfet L=3e-07 W=8e-07 AD=5.6e-14
+ AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M7@2 XI1/XI0/N2 IBRX1 VSSA_RX VSSA_RX egnfet L=3e-07 W=8e-07 AD=5.6e-14
+ AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=5.6e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M11 XI1/VBP IBRX1 VSSA_RX VSSA_RX egnfet L=3e-07 W=8e-07 AD=5.6e-14
+ AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/XI0/M11@2 XI1/VBP IBRX1 VSSA_RX VSSA_RX egnfet L=3e-07 W=8e-07 AD=5.6e-14
+ AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=5.6e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XX287/D0_noxref VSS VDDHA_TX diodenwx  AREA=2.45729e-10 perim=8.486e-05
+ sizedup=0
XX287/D1_noxref VSS VDDHA_TX diodenwx  AREA=4.01512e-10 perim=0.00035532
+ sizedup=0
XMDC2@11 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@10 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@9 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@8 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@7 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@6 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@5 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@4 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@3 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615
+ scc=0.000194942 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC2@2 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528
+ scc=0.000443878 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XX287/X22/D0_noxref VSS VDDHA_TX diodenwx  AREA=8.66626e-11 perim=5.594e-05
+ sizedup=0
XX287/X22/D1_noxref VSS XI0/XI1/N1 diodenwx  AREA=2.43222e-11 perim=2.337e-05
+ sizedup=0
XX287/X22/D2_noxref VSS VDDHA_TX diodenwx  AREA=4.32941e-10 perim=0.00010233
+ sizedup=0
XX287/X22/D3_noxref VSS VDDHA_TX diodenwx  AREA=5.235e-11 perim=2.896e-05
+ sizedup=0
XX287/X22/D4_noxref VSS XI0/XI1/XI1/XI0/N3 diodenwx  AREA=2.18474e-11
+ perim=2.022e-05 sizedup=0
XX287/X22/D5_noxref VSS VDDHA_TX diodenwx  AREA=4.89284e-10 perim=0.0001122
+ sizedup=0
XXI0/XI1/CC0 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC1 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC2 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC3 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC4 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC5 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC6 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC7 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC8 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC9 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC69 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC68 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC67 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC66 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC65 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC64 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC63 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC62 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC61 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC60 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC59 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC58 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC57 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC56 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC55 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC54 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC53 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC52 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC51 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC50 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC49 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC48 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC47 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC46 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC45 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC44 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC43 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC42 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC41 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC40 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC39 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC38 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC37 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC36 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC35 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC34 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC33 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC32 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC31 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC30 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC29 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC28 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC27 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC26 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC25 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC24 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC23 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC22 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC21 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC20 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC19 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC18 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC17 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC16 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC15 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC14 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC13 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC12 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC11 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/CC10 XI0/XI1/N1N166 XI0/VBP VSSA_TX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI1/XI1/M9 XI0/XI1/XI1/N6 XI0/XI1/XI1/N8 XI0/XI1/XI1/N1 VSSA_TX egnfet
+ L=6e-07 W=1.54e-06 AD=3.388e-13 AS=2.079e-13 PD=3.52e-06 PS=1.81e-06 M=1
+ sca=0.72776 scb=1.92596e-05 scc=1.08865e-09 lpccnr=5.55e-07 covpccnr=0
+ wrxcnr=1.386e-06 sa=2.2e-07 sb=1.09e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M9@4 XI0/XI1/XI1/N6 XI0/XI1/XI1/N8 XI0/XI1/XI1/N1 VSSA_TX egnfet
+ L=6e-07 W=1.54e-06 AD=3.388e-13 AS=2.079e-13 PD=3.52e-06 PS=1.81e-06 M=1
+ sca=0.72776 scb=1.92596e-05 scc=1.08865e-09 lpccnr=5.55e-07 covpccnr=0
+ wrxcnr=1.386e-06 sa=1.09e-06 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M9@3 XI0/XI1/XI1/N6 XI0/XI1/XI1/N8 XI0/XI1/XI1/N1 VSSA_TX egnfet
+ L=6e-07 W=1.54e-06 AD=3.388e-13 AS=2.079e-13 PD=3.52e-06 PS=1.81e-06 M=1
+ sca=0.72776 scb=1.92596e-05 scc=1.08865e-09 lpccnr=5.55e-07 covpccnr=0
+ wrxcnr=1.386e-06 sa=2.2e-07 sb=1.09e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M9@2 XI0/XI1/XI1/N6 XI0/XI1/XI1/N8 XI0/XI1/XI1/N1 VSSA_TX egnfet
+ L=6e-07 W=1.54e-06 AD=3.388e-13 AS=2.079e-13 PD=3.52e-06 PS=1.81e-06 M=1
+ sca=0.72776 scb=1.92596e-05 scc=1.08865e-09 lpccnr=5.55e-07 covpccnr=0
+ wrxcnr=1.386e-06 sa=1.09e-06 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M13 XI0/XI1/XI1/N7 XI0/XI1/PD VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=1.03966
+ scb=5.69875e-05 scc=3.99185e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M10 XI0/VBP XI0/XI1/XI1/N8 XI0/XI1/XI1/N2 VSSA_TX egnfet L=6e-07
+ W=1.54e-06 AD=3.388e-13 AS=2.079e-13 PD=3.52e-06 PS=1.81e-06 M=1 sca=0.72776
+ scb=1.92596e-05 scc=1.08865e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06
+ sa=2.2e-07 sb=1.09e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M10@4 XI0/VBP XI0/XI1/XI1/N8 XI0/XI1/XI1/N2 VSSA_TX egnfet L=6e-07
+ W=1.54e-06 AD=3.388e-13 AS=2.079e-13 PD=3.52e-06 PS=1.81e-06 M=1 sca=0.72776
+ scb=1.92596e-05 scc=1.08865e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06
+ sa=1.09e-06 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M10@3 XI0/VBP XI0/XI1/XI1/N8 XI0/XI1/XI1/N2 VSSA_TX egnfet L=6e-07
+ W=1.54e-06 AD=3.388e-13 AS=2.079e-13 PD=3.52e-06 PS=1.81e-06 M=1 sca=0.72776
+ scb=1.92596e-05 scc=1.08865e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06
+ sa=2.2e-07 sb=1.09e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M10@2 XI0/VBP XI0/XI1/XI1/N8 XI0/XI1/XI1/N2 VSSA_TX egnfet L=6e-07
+ W=1.54e-06 AD=3.388e-13 AS=2.079e-13 PD=3.52e-06 PS=1.81e-06 M=1 sca=0.72776
+ scb=1.92596e-05 scc=1.08865e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06
+ sa=1.09e-06 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M7 XI0/XI1/XI1/N6 XI0/XI1/XI1/N9 XI0/XI1/XI1/N4 VDDHA_TX egpfet
+ L=3e-07 W=3.76e-06 AD=5.076e-13 AS=8.272e-13 PD=4.03e-06 PS=7.96e-06 M=1
+ sca=2.21946 scb=0.00182982 scc=6.07933e-05 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.384e-06 sa=2.2e-07 sb=1.93e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M5 XI0/XI1/XI1/N4 XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1 sca=7.73877
+ scb=0.00749354 scc=0.000124694 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06
+ sa=2.2e-07 sb=1.93e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M7@4 XI0/XI1/XI1/N6 XI0/XI1/XI1/N9 XI0/XI1/XI1/N4 VDDHA_TX egpfet
+ L=3e-07 W=3.76e-06 AD=5.076e-13 AS=5.076e-13 PD=4.03e-06 PS=4.03e-06 M=1
+ sca=2.21946 scb=0.00182982 scc=6.07933e-05 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.384e-06 sa=7.9e-07 sb=1.36e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M5@4 XI0/XI1/XI1/N4 XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.88e-06 AD=2.538e-13 AS=2.538e-13 PD=2.15e-06 PS=2.15e-06 M=1 sca=4.26982
+ scb=0.00186931 scc=5.95167e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06
+ sa=7.9e-07 sb=1.36e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M7@3 XI0/XI1/XI1/N6 XI0/XI1/XI1/N9 XI0/XI1/XI1/N4 VDDHA_TX egpfet
+ L=3e-07 W=3.76e-06 AD=5.076e-13 AS=5.076e-13 PD=4.03e-06 PS=4.03e-06 M=1
+ sca=2.21946 scb=0.00182982 scc=6.07933e-05 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.384e-06 sa=1.36e-06 sb=7.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M5@3 XI0/XI1/XI1/N4 XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.88e-06 AD=2.538e-13 AS=2.538e-13 PD=2.15e-06 PS=2.15e-06 M=1 sca=1.32138
+ scb=0.000149054 scc=2.85087e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06
+ sa=1.36e-06 sb=7.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M7@2 XI0/XI1/XI1/N6 XI0/XI1/XI1/N9 XI0/XI1/XI1/N4 VDDHA_TX egpfet
+ L=3e-07 W=3.76e-06 AD=5.076e-13 AS=8.272e-13 PD=4.03e-06 PS=7.96e-06 M=1
+ sca=2.21946 scb=0.00182982 scc=6.07933e-05 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.384e-06 sa=1.93e-06 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/MD VDDHA_TX VDDHA_TX VDDHA_TX VDDHA_TX egpfet L=2.8e-07 W=4e-06
+ AD=8.8e-13 AS=8.8e-13 PD=8.44e-06 PS=8.44e-06 M=1 sca=2.10466 scb=0.00172003
+ scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.2e-07
+ sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M1 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet L=2.8e-07
+ W=4e-06 AD=5.4e-13 AS=8.8e-13 PD=4.27e-06 PS=8.44e-06 M=1 sca=2.10466
+ scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06
+ sa=2.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M1@16 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=7.7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M1@15 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.32e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M1@14 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.87e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M1@13 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=1.87e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M1@12 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=1.32e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M1@11 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=7.7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M1@10 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=8.8e-13 PD=4.27e-06 PS=8.44e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet L=2.8e-07
+ W=4e-06 AD=5.4e-13 AS=8.8e-13 PD=4.27e-06 PS=8.44e-06 M=1 sca=2.10466
+ scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06
+ sa=2.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2@16 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=7.7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2@15 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.32e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2@14 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.87e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2@13 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=1.87e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2@12 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=1.32e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2@11 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=7.7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2@10 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=8.8e-13 PD=4.27e-06 PS=8.44e-06 M=1
+ sca=2.10466 scb=0.00172003 scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/MD@4 VDDHA_TX VDDHA_TX VDDHA_TX VDDHA_TX egpfet L=2.8e-07 W=4e-06
+ AD=8.8e-13 AS=8.8e-13 PD=8.44e-06 PS=8.44e-06 M=1 sca=2.10466 scb=0.00172003
+ scc=5.71457e-05 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.2e-07
+ sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M8 XI0/VBP XI0/XI1/XI1/N9 XI0/XI1/XI1/N5 VDDHA_TX egpfet L=3e-07
+ W=3.76e-06 AD=5.076e-13 AS=8.272e-13 PD=4.03e-06 PS=7.96e-06 M=1 sca=2.21946
+ scb=0.00182982 scc=6.07933e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=3.384e-06
+ sa=2.2e-07 sb=1.93e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M8@4 XI0/VBP XI0/XI1/XI1/N9 XI0/XI1/XI1/N5 VDDHA_TX egpfet L=3e-07
+ W=3.76e-06 AD=5.076e-13 AS=5.076e-13 PD=4.03e-06 PS=4.03e-06 M=1 sca=2.21946
+ scb=0.00182982 scc=6.07933e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=3.384e-06
+ sa=7.9e-07 sb=1.36e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M6 XI0/XI1/XI1/N5 XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.88e-06 AD=2.538e-13 AS=2.538e-13 PD=2.15e-06 PS=2.15e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=7.9e-07 sb=1.36e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M8@3 XI0/VBP XI0/XI1/XI1/N9 XI0/XI1/XI1/N5 VDDHA_TX egpfet L=3e-07
+ W=3.76e-06 AD=5.076e-13 AS=5.076e-13 PD=4.03e-06 PS=4.03e-06 M=1 sca=2.21946
+ scb=0.00182982 scc=6.07933e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=3.384e-06
+ sa=1.36e-06 sb=7.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M6@4 XI0/XI1/XI1/N5 XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.88e-06 AD=2.538e-13 AS=2.538e-13 PD=2.15e-06 PS=2.15e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.36e-06 sb=7.9e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M8@2 XI0/VBP XI0/XI1/XI1/N9 XI0/XI1/XI1/N5 VDDHA_TX egpfet L=3e-07
+ W=3.76e-06 AD=5.076e-13 AS=8.272e-13 PD=4.03e-06 PS=7.96e-06 M=1 sca=2.21946
+ scb=0.00182982 scc=6.07933e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=3.384e-06
+ sa=1.93e-06 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M6@3 XI0/XI1/XI1/N5 XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.93e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX287/X22/X117/D0_noxref VSS VDDHA_TX diodenwx  AREA=4.87035e-11 perim=2.792e-05
+ sizedup=0
XXI0/XI1/RRC1 XI0/XI1/N1N166 X287/X22/X117/noxref_11 VDDHA_TX opppcres 2452.51
+ M=1 w=2e-06 l=8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/RRC2 XI0/XI1/N1N69 X287/X22/X117/noxref_11 VDDHA_TX opppcres 2452.51
+ M=1 w=2e-06 l=8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/RRTMP XI0/FB XI0/XI1/N1N69 VSSA_TX opppcres 772.179 M=1 w=2e-06
+ l=2.43e-06   bp=3 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/M2 XI0/FB IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=1.53e-13 PD=1.12e-06 PS=2.14e-06 M=1 sca=0.865276 scb=3.01673e-05
+ scc=1.66086e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=1.7e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M2@8 XI0/FB IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=1.53e-13 PD=1.12e-06 PS=2.14e-06 M=1 sca=0.600443 scb=2.85471e-05
+ scc=2.43563e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=1.7e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M2@7 XI0/FB IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.865276 scb=3.01673e-05
+ scc=1.66086e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=7.9e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M2@6 XI0/FB IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.941871 scb=4.47798e-05
+ scc=3.82059e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=7.9e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M2@5 XI0/FB IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.865276 scb=3.01673e-05
+ scc=1.66086e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=1.41e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M2@4 XI0/FB IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.941871 scb=4.47798e-05
+ scc=3.82059e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=1.41e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M2@3 XI0/FB IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.865276 scb=3.01673e-05
+ scc=1.66086e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M2@2 XI0/FB IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.941871 scb=4.47798e-05
+ scc=3.82059e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M0 IBTX2 IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.865276 scb=3.01673e-05
+ scc=1.66086e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M0@8 IBTX2 IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.941871 scb=4.47798e-05
+ scc=3.82059e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M0@7 IBTX2 IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.865276 scb=3.01673e-05
+ scc=1.66086e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06
+ sb=1.41e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M0@6 IBTX2 IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.941871 scb=4.47798e-05
+ scc=3.82059e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06
+ sb=1.41e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M0@5 IBTX2 IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.865276 scb=3.01673e-05
+ scc=1.66086e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06
+ sb=7.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M0@4 IBTX2 IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=9.9e-14 PD=1.12e-06 PS=1.12e-06 M=1 sca=0.941871 scb=4.47798e-05
+ scc=3.82059e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06
+ sb=7.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M0@3 IBTX2 IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=1.53e-13 PD=1.12e-06 PS=2.14e-06 M=1 sca=0.865276 scb=3.01673e-05
+ scc=1.66086e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06
+ sb=1.7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M0@2 IBTX2 IBTX2 VSSA_TX VSSA_TX egnfet L=4e-07 W=9e-07 AD=9.9e-14
+ AS=1.53e-13 PD=1.12e-06 PS=2.14e-06 M=1 sca=0.941871 scb=4.47798e-05
+ scc=3.82059e-09 lpccnr=3.75e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06
+ sb=1.7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M4 IBTX2 XI0/XI1/PD VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=6.8e-14
+ AS=6.8e-14 PD=1.14e-06 PS=1.14e-06 M=1 sca=1.12547 scb=8.00455e-05
+ scc=8.19324e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.7e-07 sb=1.7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M3 XI0/XI1/N1N69 VSSA_TX XI0/XI1/N1 XI0/XI1/N1 egpfet L=1.5e-07
+ W=7.56e-06 AD=8.316e-13 AS=1.2852e-12 PD=7.78e-06 PS=1.546e-05 M=1 sca=9.37165
+ scb=0.00719944 scc=8.50181e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=6.804e-06
+ sa=1.7e-07 sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M3@2 XI0/XI1/N1N69 VSSA_TX XI0/XI1/N1 XI0/XI1/N1 egpfet L=1.5e-07
+ W=7.56e-06 AD=8.316e-13 AS=1.2852e-12 PD=7.78e-06 PS=1.546e-05 M=1 sca=9.37165
+ scb=0.00719944 scc=8.50181e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=6.804e-06
+ sa=5.4e-07 sb=1.7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M1 XI0/XI1/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07 W=5e-06
+ AD=5.5e-13 AS=8.5e-13 PD=5.22e-06 PS=1.034e-05 M=1 sca=6.96176 scb=0.00571125
+ scc=7.06854e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.7e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M1@10 XI0/XI1/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07 W=5e-06
+ AD=5.5e-13 AS=5.5e-13 PD=5.22e-06 PS=5.22e-06 M=1 sca=4.57898 scb=0.00214689
+ scc=2.67197e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=6.9e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M1@9 XI0/XI1/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07 W=5e-06
+ AD=5.5e-13 AS=5.5e-13 PD=5.22e-06 PS=5.22e-06 M=1 sca=3.67336 scb=0.00148648
+ scc=2.5714e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.21e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M1@8 XI0/XI1/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07 W=5e-06
+ AD=5.5e-13 AS=5.5e-13 PD=5.22e-06 PS=5.22e-06 M=1 sca=2.39938 scb=0.00135711
+ scc=2.56929e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.73e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M1@7 XI0/XI1/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07 W=5e-06
+ AD=5.5e-13 AS=5.5e-13 PD=5.22e-06 PS=5.22e-06 M=1 sca=2.39938 scb=0.00135711
+ scc=2.56929e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M1@6 XI0/XI1/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07 W=5e-06
+ AD=5.5e-13 AS=5.5e-13 PD=5.22e-06 PS=5.22e-06 M=1 sca=2.39938 scb=0.00135711
+ scc=2.56929e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M1@5 XI0/XI1/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07 W=5e-06
+ AD=5.5e-13 AS=5.5e-13 PD=5.22e-06 PS=5.22e-06 M=1 sca=2.39938 scb=0.00135711
+ scc=2.56929e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.73e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M1@4 XI0/XI1/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07 W=5e-06
+ AD=5.5e-13 AS=5.5e-13 PD=5.22e-06 PS=5.22e-06 M=1 sca=3.59633 scb=0.00145801
+ scc=2.57053e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.21e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M1@3 XI0/XI1/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07 W=5e-06
+ AD=5.5e-13 AS=5.5e-13 PD=5.22e-06 PS=5.22e-06 M=1 sca=4.40877 scb=0.00197902
+ scc=2.63044e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=6.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M1@2 XI0/XI1/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07 W=5e-06
+ AD=5.5e-13 AS=8.5e-13 PD=5.22e-06 PS=1.034e-05 M=1 sca=6.45782 scb=0.00484809
+ scc=5.2992e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/RRD1 VDDHA_TX VDDHA_TX VDDHA_TX opppcres 4877.98 M=1 w=1e-06
+ l=7.91e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/XI1/RR1 X287/X22/X118/noxref_13 VSSA_TX VDDHA_TX opppcres 1034.64
+ M=1 w=2e-06 l=3.3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/RR1 IBTX1 XI0/XI1/XI0/VCM7 VDDHA_TX opppcres 944.134 M=1 w=2e-06
+ l=3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/XI1/RR2 X287/X22/X118/noxref_13 X287/X22/X118/noxref_14 VDDHA_TX
+ opppcres 1034.64 M=1 w=2e-06 l=3.3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/RR2 XI0/XI1/XI0/VCM6 XI0/XI1/XI0/VCM7 VDDHA_TX opppcres 944.134 M=1
+ w=2e-06 l=3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/XI1/RR3 X287/X22/X118/noxref_15 X287/X22/X118/noxref_14 VDDHA_TX
+ opppcres 1034.64 M=1 w=2e-06 l=3.3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/RR3 XI0/XI1/XI0/VCM6 XI0/XI1/XI0/VCM5 VDDHA_TX opppcres 944.134 M=1
+ w=2e-06 l=3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/XI1/RR4 X287/X22/X118/noxref_15 X287/X22/X118/noxref_16 VDDHA_TX
+ opppcres 1034.64 M=1 w=2e-06 l=3.3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/RR4 XI0/XI1/XI0/VCM4 XI0/XI1/XI0/VCM5 VDDHA_TX opppcres 944.134 M=1
+ w=2e-06 l=3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/XI1/RR5 X287/X22/X118/noxref_17 X287/X22/X118/noxref_16 VDDHA_TX
+ opppcres 1034.64 M=1 w=2e-06 l=3.3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/RR5 XI0/XI1/XI0/VCM4 XI0/XI1/XI0/VCM3 VDDHA_TX opppcres 944.134 M=1
+ w=2e-06 l=3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/XI1/RR6 X287/X22/X118/noxref_17 X287/X22/X118/noxref_18 VDDHA_TX
+ opppcres 1034.64 M=1 w=2e-06 l=3.3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/RR6 XI0/XI1/XI0/VCM2 XI0/XI1/XI0/VCM3 VDDHA_TX opppcres 944.134 M=1
+ w=2e-06 l=3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/XI1/RR7 X287/X22/X118/noxref_19 X287/X22/X118/noxref_18 VDDHA_TX
+ opppcres 1034.64 M=1 w=2e-06 l=3.3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/RR7 XI0/XI1/XI0/VCM2 XI0/XI1/XI0/VCM1 VDDHA_TX opppcres 944.134 M=1
+ w=2e-06 l=3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/XI1/RR8 X287/X22/X118/noxref_19 XI0/XI1/XI0/VCM0 VDDHA_TX opppcres
+ 1034.64 M=1 w=2e-06 l=3.3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/RR8 XI0/XI1/XI0/VCM0 XI0/XI1/XI0/VCM1 VDDHA_TX opppcres 944.134 M=1
+ w=2e-06 l=3e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/RRD3 VDDHA_TX VDDHA_TX VDDHA_TX opppcres 15338.2 M=1 w=1e-06
+ l=2.515e-05   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/RRD4 VDDHA_TX VDDHA_TX VDDHA_TX opppcres 15338.2 M=1 w=1e-06
+ l=2.515e-05   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/XI0/RRD2 VDDHA_TX VDDHA_TX VDDHA_TX opppcres 4877.98 M=1 w=1e-06
+ l=7.91e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI1/M19C VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@36 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@35 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@34 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@33 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@32 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@31 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@30 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@29 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@28 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@27 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@26 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@25 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@24 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@23 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@22 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@32 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@31 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@30 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@29 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@28 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@27 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@26 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@25 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@24 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@23 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@22 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@21 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@20 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@19 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@18 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19A VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@48 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@47 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@46 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@45 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@44 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@43 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@42 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@41 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@40 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@39 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@38 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@37 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@36 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@35 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@34 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@33 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@32 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@31 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@30 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@29 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@28 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@27 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@26 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0.608318 scb=6.93782e-05
+ scc=6.17333e-08 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@21 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@20 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@19 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@18 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@17 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@16 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@15 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@14 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@13 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@12 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@11 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@10 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@9 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@8 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@7 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@6 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@17 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@5 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@16 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@4 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@15 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@14 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@13 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@12 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@11 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@10 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@9 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@8 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@7 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@6 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@5 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@4 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@3 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@3 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=3.5e-13
+ AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19B@2 VSSA_TX IBTX1 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19C@2 VSSA_TX IBTX2 VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@25 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@24 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@23 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@22 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@21 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@20 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@19 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@18 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/M19A@17 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@16 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@15 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@14 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@13 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@12 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@11 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@10 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@9 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@8 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@7 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@6 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@5 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@4 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@3 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M19A@2 VSSA_TX XI0/VCM VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.86012 scb=0.00154221
+ scc=5.96657e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M18 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=6.62202 scb=0.005221
+ scc=0.000567173 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M18@2 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@3 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=4.7619 scb=0.00367879
+ scc=0.000507507 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M18@4 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@5 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@6 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@7 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@8 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@9 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@10 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@11 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@12 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@13 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@14 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@15 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@16 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@17 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=4.7619 scb=0.00367879
+ scc=0.000507507 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M18@18 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@19 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=4.7619 scb=0.00367879
+ scc=0.000507507 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M18@20 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=4.06065 scb=0.00349225
+ scc=0.000163631 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M18@21 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.86012 scb=0.00154221
+ scc=5.96657e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M18@22 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M18@23 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@24 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M18@25 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@26 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M18@27 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@28 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/M18@29 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M18@30 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@2 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/MC1@3 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@4 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/MC1@5 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@6 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/MC1@7 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@8 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/MC1@9 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@10 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/MC1@11 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@12 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/MC1@13 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@14 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/MC1@15 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@16 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/MC1@17 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@18 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/MC1@19 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.20053 scb=0.00195005
+ scc=0.000103965 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@20 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/MC1@21 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=2.29354 scb=0.00202716
+ scc=0.000106948 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@22 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX287/X22/X120/D0_noxref VSS VDDHA_TX diodenwx  AREA=7.6725e-11 perim=4.842e-05
+ sizedup=0
XXI0/XI1/XI0/XI0/XG0/M2 XI0/XI1/XI0/XI0/N1N140 XI0/CCMH0 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI0/XI0/XG2/M2 XI0/XI1/XI0/XI0/N1N134 XI0/CCMH1 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI0/XI0/XG1/M2 XI0/XI1/XI0/XI0/COI XI0/XI1/XI0/XI0/N1N140 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06
+ M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XG3/M2 XI0/XI1/XI0/XI0/C1I XI0/XI1/XI0/XI0/N1N134 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06
+ M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XG4/M2 XI0/XI1/XI0/XI0/SHB XI0/CCMH2 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/MHN XI0/XI1/XI0/XI0/N1 XI0/XI1/XI0/XI0/SH XI0/VCM VSSA_TX
+ egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/M3N XI0/XI1/XI0/VCM7 XI0/XI1/XI0/XI0/XI1/S3
+ XI0/XI1/XI0/XI0/N1 VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG11/M2 XI0/XI1/XI0/XI0/XI1/S3B XI0/XI1/XI0/XI0/XI1/S3
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/M2N XI0/XI1/XI0/VCM6 XI0/XI1/XI0/XI0/XI1/S2
+ XI0/XI1/XI0/XI0/N1 VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG8/M2 XI0/XI1/XI0/XI0/XI1/S2B XI0/XI1/XI0/XI0/XI1/S2
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/M1N XI0/XI1/XI0/VCM5 XI0/XI1/XI0/XI0/XI1/S1
+ XI0/XI1/XI0/XI0/N1 VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG5/M2 XI0/XI1/XI0/XI0/XI1/S1B XI0/XI1/XI0/XI0/XI1/S1
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/M0N XI0/XI1/XI0/VCM4 XI0/XI1/XI0/XI0/XI1/S0
+ XI0/XI1/XI0/XI0/N1 VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG2/M2 XI0/XI1/XI0/XI0/XI1/S0 XI0/XI1/XI0/XI0/XI1/S0B
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XG5/M2 XI0/XI1/XI0/XI0/SH XI0/XI1/XI0/XI0/SHB VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/MLN XI0/XI1/XI0/XI0/N2 XI0/XI1/XI0/XI0/SHB XI0/VCM VSSA_TX
+ egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/M3N XI0/XI1/XI0/VCM3 XI0/XI1/XI0/XI0/XI0/S3
+ XI0/XI1/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG11/M2 XI0/XI1/XI0/XI0/XI0/S3B XI0/XI1/XI0/XI0/XI0/S3
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/M2N XI0/XI1/XI0/VCM2 XI0/XI1/XI0/XI0/XI0/S2
+ XI0/XI1/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG8/M2 XI0/XI1/XI0/XI0/XI0/S2B XI0/XI1/XI0/XI0/XI0/S2
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/M1N XI0/XI1/XI0/VCM1 XI0/XI1/XI0/XI0/XI0/S1
+ XI0/XI1/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG5/M2 XI0/XI1/XI0/XI0/XI0/S1B XI0/XI1/XI0/XI0/XI0/S1
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/M0N XI0/XI1/XI0/VCM0 XI0/XI1/XI0/XI0/XI0/S0
+ XI0/XI1/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG2/M2 XI0/XI1/XI0/XI0/XI0/S0 XI0/XI1/XI0/XI0/XI0/S0B
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XG0/M1 XI0/XI1/XI0/XI0/N1N140 XI0/CCMH0 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1
+ sca=9.87748 scb=0.00793829 scc=0.000299729 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XG2/M1 XI0/XI1/XI0/XI0/N1N134 XI0/CCMH1 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1
+ sca=8.3546 scb=0.0065938 scc=0.000296143 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XG1/M1 XI0/XI1/XI0/XI0/COI XI0/XI1/XI0/XI0/N1N140 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06
+ PS=3.04e-06 M=1 sca=7.12959 scb=0.00648536 scc=0.000296129 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XG3/M1 XI0/XI1/XI0/XI0/C1I XI0/XI1/XI0/XI0/N1N134 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06
+ PS=3.04e-06 M=1 sca=7.12959 scb=0.00648536 scc=0.000296129 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG9/M2 XI0/XI1/XI0/XI0/XI1/N4 XI0/XI1/XI0/XI0/COI VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06
+ PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG9/M1 XI0/XI1/XI0/XI0/XI1/N4 XI0/XI1/XI0/XI0/C1I VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06
+ PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.26e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XG4/M1 XI0/XI1/XI0/XI0/SHB XI0/CCMH2 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1
+ sca=6.51926 scb=0.00389739 scc=7.76568e-05 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG10/M1 XI0/XI1/XI0/XI0/XI1/S3 XI0/XI1/XI0/XI0/XI1/N4
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG13/M1 XI0/XI1/XI0/XI0/XI1/C0B XI0/XI1/XI0/XI0/COI
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG4/M1 XI0/XI1/XI0/XI0/XI1/S1 XI0/XI1/XI0/XI0/XI1/N2
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG5/M1 XI0/XI1/XI0/XI0/XI1/S1B XI0/XI1/XI0/XI0/XI1/S1
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=5.17805 scb=0.00374279 scc=7.76283e-05
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG0/M1 XI0/XI1/XI0/XI0/XI1/XG0/N1 XI0/XI1/XI0/XI0/COI
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13
+ PD=1.54e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/M0P XI0/XI1/XI0/VCM4 XI0/XI1/XI0/XI0/XI1/S0B
+ XI0/XI1/XI0/XI0/N1 VDDHA_TX egpfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=7.24638 scb=0.00892862 scc=0.00025501
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG0/M2 XI0/XI1/XI0/XI0/XI1/N1 XI0/XI1/XI0/XI0/C1I
+ XI0/XI1/XI0/XI0/XI1/XG0/N1 VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13
+ AS=9.8e-14 PD=3.04e-06 PS=1.54e-06 M=1 sca=7.25571 scb=0.00665164
+ scc=0.000316017 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=4.1e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG2/M1 XI0/XI1/XI0/XI0/XI1/S0 XI0/XI1/XI0/XI0/XI1/S0B
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=5.17805 scb=0.00374279 scc=7.76283e-05
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG1/M1 XI0/XI1/XI0/XI0/XI1/S0B XI0/XI1/XI0/XI0/XI1/N1
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG9/M2 XI0/XI1/XI0/XI0/XI0/N4 XI0/XI1/XI0/XI0/COI VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06
+ PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG9/M1 XI0/XI1/XI0/XI0/XI0/N4 XI0/XI1/XI0/XI0/C1I VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06
+ PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.26e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XG5/M1 XI0/XI1/XI0/XI0/SH XI0/XI1/XI0/XI0/SHB VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1
+ sca=5.17805 scb=0.00374279 scc=7.76283e-05 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG10/M1 XI0/XI1/XI0/XI0/XI0/S3 XI0/XI1/XI0/XI0/XI0/N4
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG13/M1 XI0/XI1/XI0/XI0/XI0/C0B XI0/XI1/XI0/XI0/COI
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG4/M1 XI0/XI1/XI0/XI0/XI0/S1 XI0/XI1/XI0/XI0/XI0/N2
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG5/M1 XI0/XI1/XI0/XI0/XI0/S1B XI0/XI1/XI0/XI0/XI0/S1
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=5.17805 scb=0.00374279 scc=7.76283e-05
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG0/M1 XI0/XI1/XI0/XI0/XI0/XG0/N1 XI0/XI1/XI0/XI0/COI
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13
+ PD=1.54e-06 PS=3.04e-06 M=1 sca=8.78954 scb=0.00690469 scc=0.000316098
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/M0P XI0/XI1/XI0/VCM0 XI0/XI1/XI0/XI0/XI0/S0B
+ XI0/XI1/XI0/XI0/N2 VDDHA_TX egpfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=8.78784 scb=0.00918614 scc=0.000255095
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG0/M2 XI0/XI1/XI0/XI0/XI0/N1 XI0/XI1/XI0/XI0/C1I
+ XI0/XI1/XI0/XI0/XI0/XG0/N1 VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13
+ AS=9.8e-14 PD=3.04e-06 PS=1.54e-06 M=1 sca=9.34792 scb=0.00734253
+ scc=0.000316727 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=4.1e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG2/M1 XI0/XI1/XI0/XI0/XI0/S0 XI0/XI1/XI0/XI0/XI0/S0B
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=9.09753 scb=0.00698282 scc=9.89973e-05
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG1/M1 XI0/XI1/XI0/XI0/XI0/S0B XI0/XI1/XI0/XI0/XI0/N1
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=15.3855 scb=0.017138 scc=0.000637805
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/MHP XI0/XI1/XI0/XI0/N1 XI0/XI1/XI0/XI0/SHB XI0/VCM VDDHA_TX
+ egpfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=7.24638 scb=0.00892862 scc=0.00025501 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG9/M4 XI0/XI1/XI0/XI0/XI1/XG9/N1 XI0/XI1/XI0/XI0/COI
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07
+ PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG9/M3 XI0/XI1/XI0/XI0/XI1/N4 XI0/XI1/XI0/XI0/C1I
+ XI0/XI1/XI0/XI0/XI1/XG9/N1 VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=9.6e-14
+ AS=5.6e-14 PD=1.84e-06 PS=9.4e-07 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG10/M2 XI0/XI1/XI0/XI0/XI1/S3 XI0/XI1/XI0/XI0/XI1/N4
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG13/M2 XI0/XI1/XI0/XI0/XI1/C0B XI0/XI1/XI0/XI0/COI VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06
+ M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG6/M4 XI0/XI1/XI0/XI0/XI1/XG6/N1 XI0/XI1/XI0/XI0/XI1/C0B
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07
+ PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG6/M3 XI0/XI1/XI0/XI0/XI1/N3 XI0/XI1/XI0/XI0/C1I
+ XI0/XI1/XI0/XI0/XI1/XG6/N1 VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=9.6e-14
+ AS=5.6e-14 PD=1.84e-06 PS=9.4e-07 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG7/M2 XI0/XI1/XI0/XI0/XI1/S2 XI0/XI1/XI0/XI0/XI1/N3
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG12/M2 XI0/XI1/XI0/XI0/XI1/C1B XI0/XI1/XI0/XI0/C1I VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06
+ M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG3/M4 XI0/XI1/XI0/XI0/XI1/XG3/N1 XI0/XI1/XI0/XI0/COI
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07
+ PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG3/M3 XI0/XI1/XI0/XI0/XI1/N2 XI0/XI1/XI0/XI0/XI1/C1B
+ XI0/XI1/XI0/XI0/XI1/XG3/N1 VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=9.6e-14
+ AS=5.6e-14 PD=1.84e-06 PS=9.4e-07 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG4/M2 XI0/XI1/XI0/XI0/XI1/S1 XI0/XI1/XI0/XI0/XI1/N2
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG0/M3 XI0/XI1/XI0/XI0/XI1/N1 XI0/XI1/XI0/XI0/COI VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06
+ M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG0/M4 XI0/XI1/XI0/XI0/XI1/N1 XI0/XI1/XI0/XI0/C1I VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06
+ M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=4.1e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG1/M2 XI0/XI1/XI0/XI0/XI1/S0B XI0/XI1/XI0/XI0/XI1/N1
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG6/M2 XI0/XI1/XI0/XI0/XI1/N3 XI0/XI1/XI0/XI0/XI1/C0B
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13
+ PD=1.54e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/M3P XI0/XI1/XI0/VCM7 XI0/XI1/XI0/XI0/XI1/S3B
+ XI0/XI1/XI0/XI0/N1 VDDHA_TX egpfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=7.24638 scb=0.00892862 scc=0.00025501
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG6/M1 XI0/XI1/XI0/XI0/XI1/N3 XI0/XI1/XI0/XI0/C1I VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06
+ PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.26e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG11/M1 XI0/XI1/XI0/XI0/XI1/S3B XI0/XI1/XI0/XI0/XI1/S3
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=5.17805 scb=0.00374279 scc=7.76283e-05
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG7/M1 XI0/XI1/XI0/XI0/XI1/S2 XI0/XI1/XI0/XI0/XI1/N3
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/M2P XI0/XI1/XI0/VCM6 XI0/XI1/XI0/XI0/XI1/S2B
+ XI0/XI1/XI0/XI0/N1 VDDHA_TX egpfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=7.24638 scb=0.00892862 scc=0.00025501
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG12/M1 XI0/XI1/XI0/XI0/XI1/C1B XI0/XI1/XI0/XI0/C1I
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG8/M1 XI0/XI1/XI0/XI0/XI1/S2B XI0/XI1/XI0/XI0/XI1/S2
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=5.17805 scb=0.00374279 scc=7.76283e-05
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG3/M2 XI0/XI1/XI0/XI0/XI1/N2 XI0/XI1/XI0/XI0/COI VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06
+ PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/XG3/M1 XI0/XI1/XI0/XI0/XI1/N2 XI0/XI1/XI0/XI0/XI1/C1B
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13
+ PD=1.54e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI1/M1P XI0/XI1/XI0/VCM5 XI0/XI1/XI0/XI0/XI1/S1B
+ XI0/XI1/XI0/XI0/N1 VDDHA_TX egpfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=7.24638 scb=0.00892862 scc=0.00025501
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/MLP XI0/XI1/XI0/XI0/N2 XI0/XI1/XI0/XI0/SH XI0/VCM VDDHA_TX
+ egpfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=7.24638 scb=0.00892862 scc=0.00025501 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG9/M4 XI0/XI1/XI0/XI0/XI0/XG9/N1 XI0/XI1/XI0/XI0/COI
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07
+ PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG9/M3 XI0/XI1/XI0/XI0/XI0/N4 XI0/XI1/XI0/XI0/C1I
+ XI0/XI1/XI0/XI0/XI0/XG9/N1 VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=9.6e-14
+ AS=5.6e-14 PD=1.84e-06 PS=9.4e-07 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG10/M2 XI0/XI1/XI0/XI0/XI0/S3 XI0/XI1/XI0/XI0/XI0/N4
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG13/M2 XI0/XI1/XI0/XI0/XI0/C0B XI0/XI1/XI0/XI0/COI VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06
+ M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG6/M4 XI0/XI1/XI0/XI0/XI0/XG6/N1 XI0/XI1/XI0/XI0/XI0/C0B
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07
+ PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG6/M3 XI0/XI1/XI0/XI0/XI0/N3 XI0/XI1/XI0/XI0/C1I
+ XI0/XI1/XI0/XI0/XI0/XG6/N1 VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=9.6e-14
+ AS=5.6e-14 PD=1.84e-06 PS=9.4e-07 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG7/M2 XI0/XI1/XI0/XI0/XI0/S2 XI0/XI1/XI0/XI0/XI0/N3
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG12/M2 XI0/XI1/XI0/XI0/XI0/C1B XI0/XI1/XI0/XI0/C1I VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06
+ M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG3/M4 XI0/XI1/XI0/XI0/XI0/XG3/N1 XI0/XI1/XI0/XI0/COI
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07
+ PS=1.84e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG3/M3 XI0/XI1/XI0/XI0/XI0/N2 XI0/XI1/XI0/XI0/XI0/C1B
+ XI0/XI1/XI0/XI0/XI0/XG3/N1 VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=9.6e-14
+ AS=5.6e-14 PD=1.84e-06 PS=9.4e-07 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG4/M2 XI0/XI1/XI0/XI0/XI0/S1 XI0/XI1/XI0/XI0/XI0/N2
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG0/M3 XI0/XI1/XI0/XI0/XI0/N1 XI0/XI1/XI0/XI0/COI VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06
+ M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG0/M4 XI0/XI1/XI0/XI0/XI0/N1 XI0/XI1/XI0/XI0/C1I VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06
+ M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=4.1e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG1/M2 XI0/XI1/XI0/XI0/XI0/S0B XI0/XI1/XI0/XI0/XI0/N1
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG6/M2 XI0/XI1/XI0/XI0/XI0/N3 XI0/XI1/XI0/XI0/XI0/C0B
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13
+ PD=1.54e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/M3P XI0/XI1/XI0/VCM3 XI0/XI1/XI0/XI0/XI0/S3B
+ XI0/XI1/XI0/XI0/N2 VDDHA_TX egpfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=7.24638 scb=0.00892862 scc=0.00025501
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG6/M1 XI0/XI1/XI0/XI0/XI0/N3 XI0/XI1/XI0/XI0/C1I VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06
+ PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.26e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG11/M1 XI0/XI1/XI0/XI0/XI0/S3B XI0/XI1/XI0/XI0/XI0/S3
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=5.17805 scb=0.00374279 scc=7.76283e-05
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG7/M1 XI0/XI1/XI0/XI0/XI0/S2 XI0/XI1/XI0/XI0/XI0/N3
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/M2P XI0/XI1/XI0/VCM2 XI0/XI1/XI0/XI0/XI0/S2B
+ XI0/XI1/XI0/XI0/N2 VDDHA_TX egpfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=7.24638 scb=0.00892862 scc=0.00025501
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG12/M1 XI0/XI1/XI0/XI0/XI0/C1B XI0/XI1/XI0/XI0/C1I
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG8/M1 XI0/XI1/XI0/XI0/XI0/S2B XI0/XI1/XI0/XI0/XI0/S2
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13
+ PD=3.04e-06 PS=3.04e-06 M=1 sca=5.17805 scb=0.00374279 scc=7.76283e-05
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG3/M2 XI0/XI1/XI0/XI0/XI0/N2 XI0/XI1/XI0/XI0/COI VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06
+ PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/XG3/M1 XI0/XI1/XI0/XI0/XI0/N2 XI0/XI1/XI0/XI0/XI0/C1B
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13
+ PD=1.54e-06 PS=3.04e-06 M=1 sca=7.25571 scb=0.00665164 scc=0.000316017
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI0/XI0/XI0/M1P XI0/XI1/XI0/VCM1 XI0/XI1/XI0/XI0/XI0/S1B
+ XI0/XI1/XI0/XI0/N2 VDDHA_TX egpfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14
+ PD=1.04e-06 PS=1.04e-06 M=1 sca=7.24638 scb=0.00892862 scc=0.00025501
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/M6 XI0/XI1/XI1/N14 XI0/XI1/PD VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/M7 XI0/XI1/XI1/XI0/N4 XI0/XI1/PD VSSA_TX VSSA_TX egnfet
+ L=4.2e-07 W=2.5e-06 AD=3.4005e-13 AS=5.551e-13 PD=2.8e-06 PS=5.5e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=3.93e-07 covpccnr=0 wrxcnr=2.25003e-06 sa=2.2e-07
+ sb=9.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/M8 XI0/XI1/XI1/XI0/N4 XI0/XI1/XI1/N14 VSSA_TX VSSA_TX egnfet
+ L=4.2e-07 W=2.5e-06 AD=3.4005e-13 AS=5.551e-13 PD=2.8e-06 PS=5.5e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=3.93e-07 covpccnr=0 wrxcnr=2.25003e-06 sa=9.1e-07
+ sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/M1 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/N14 VSSA_TX VSSA_TX egnfet
+ L=7e-07 W=4.6e-07 AD=6.21e-14 AS=1.012e-13 PD=7.3e-07 PS=1.36e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=2.2e-07 sb=1.19e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M1@2 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/N14 VSSA_TX VSSA_TX egnfet
+ L=7e-07 W=4.6e-07 AD=6.21e-14 AS=1.012e-13 PD=7.3e-07 PS=1.36e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=1.19e-06 sb=2.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M5 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/XI0/N4 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/X1I44/M0 XI0/XI1/XI1/XI0/TIEL XI0/XI1/XI1/XI0/X1I44/N1N50
+ VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/M2 XI0/XI1/XI1/N14 XI0/XI1/XI1/N14 VSSA_TX VSSA_TX egnfet
+ L=7e-07 W=4.6e-07 AD=6.21e-14 AS=1.012e-13 PD=7.3e-07 PS=1.36e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=2.2e-07 sb=1.19e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M2@2 XI0/XI1/XI1/N14 XI0/XI1/XI1/N14 VSSA_TX VSSA_TX egnfet
+ L=7e-07 W=4.6e-07 AD=6.21e-14 AS=1.012e-13 PD=7.3e-07 PS=1.36e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=1.19e-06 sb=2.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M10 XI0/XI1/XI1/XI0/N4 XI0/XI1/XI1/N14 XI0/XI1/XI1/XI0/N1N5
+ VDDHA_TX egpfet L=2.5e-06 W=4.2e-07 AD=9.92e-14 AS=9.92e-14 PD=1.36e-06
+ PS=1.36e-06 M=1 sca=23.4834 scb=0.0244359 scc=0.00287516 lpccnr=2.265e-06
+ covpccnr=0 wrxcnr=3.78007e-07 sa=2.2e-07 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/M10@2 XI0/XI1/XI1/XI0/N4 XI0/XI1/XI1/N14 XI0/XI1/XI1/XI0/N1N5
+ VDDHA_TX egpfet L=2.5e-06 W=4.2e-07 AD=9.92e-14 AS=9.92e-14 PD=1.36e-06
+ PS=1.36e-06 M=1 sca=6.21744 scb=0.00494713 scc=4.9798e-05 lpccnr=2.265e-06
+ covpccnr=0 wrxcnr=3.78007e-07 sa=2.2e-07 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/M9 XI0/XI1/XI1/XI0/N1N5 XI0/XI1/PD VDDHA_TX VDDHA_TX egpfet
+ L=2.5e-06 W=4.2e-07 AD=9.92e-14 AS=9.92e-14 PD=1.36e-06 PS=1.36e-06 M=1
+ sca=3.22278 scb=0.00141699 scc=1.76183e-05 lpccnr=2.265e-06 covpccnr=0
+ wrxcnr=3.78007e-07 sa=2.2e-07 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/M9@2 XI0/XI1/XI1/XI0/N1N5 XI0/XI1/PD VDDHA_TX VDDHA_TX egpfet
+ L=2.5e-06 W=4.2e-07 AD=9.92e-14 AS=9.92e-14 PD=1.36e-06 PS=1.36e-06 M=1
+ sca=2.10126 scb=0.0013377 scc=1.76101e-05 lpccnr=2.265e-06 covpccnr=0
+ wrxcnr=3.78007e-07 sa=2.2e-07 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/MR XI0/XI1/XI1/XI0/N3 XI0/XI1/XI1/XI0/TIEL VDDHA_TX VDDHA_TX
+ egpfet L=8e-07 W=5.2e-07 AD=1.144e-13 AS=1.144e-13 PD=1.48e-06 PS=1.48e-06 M=1
+ sca=0 scb=0 scc=0 lpccnr=7.35e-07 covpccnr=0 wrxcnr=4.68e-07 sa=2.2e-07
+ sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/M3 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/XI0/N2 VDDHA_TX VDDHA_TX
+ egpfet L=5.4e-07 W=1.2e-06 AD=1.62e-13 AS=2.64e-13 PD=1.47e-06 PS=2.84e-06 M=1
+ sca=10.7592 scb=0.0114771 scc=0.00106852 lpccnr=5.01e-07 covpccnr=0
+ wrxcnr=1.08e-06 sa=2.2e-07 sb=1.03e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/M3@2 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/XI0/N2 VDDHA_TX VDDHA_TX
+ egpfet L=5.4e-07 W=1.2e-06 AD=1.62e-13 AS=2.64e-13 PD=1.47e-06 PS=2.84e-06 M=1
+ sca=12.2802 scb=0.0117414 scc=0.00106864 lpccnr=5.01e-07 covpccnr=0
+ wrxcnr=1.08e-06 sa=1.03e-06 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/XI0/X1I44/M1 XI0/XI1/XI1/XI0/X1I44/N1N50
+ XI0/XI1/XI1/XI0/X1I44/N1N50 VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=59.4525 scb=0.0550273
+ scc=0.00911315 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M4 XI0/XI1/XI1/N14 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/XI0/N3
+ XI0/XI1/XI1/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=1.62e-13 AS=2.64e-13
+ PD=1.47e-06 PS=2.84e-06 M=1 sca=17.3113 scb=0.0168035 scc=0.00114318
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.2e-07 sb=1.03e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M4@8 XI0/XI1/XI1/N14 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/XI0/N3
+ XI0/XI1/XI1/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=1.62e-13 AS=2.64e-13
+ PD=1.47e-06 PS=2.84e-06 M=1 sca=7.68921 scb=0.0054437 scc=7.47049e-05
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.2e-07 sb=1.03e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M4@7 XI0/XI1/XI1/N14 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/XI0/N3
+ XI0/XI1/XI1/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=1.62e-13 AS=2.64e-13
+ PD=1.47e-06 PS=2.84e-06 M=1 sca=6.5521 scb=0.00532637 scc=7.46664e-05
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.2e-07 sb=1.03e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M4@6 XI0/XI1/XI1/N14 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/XI0/N3
+ XI0/XI1/XI1/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=1.62e-13 AS=2.64e-13
+ PD=1.47e-06 PS=2.84e-06 M=1 sca=9.16105 scb=0.00687439 scc=8.49142e-05
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.2e-07 sb=1.03e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M4@5 XI0/XI1/XI1/N14 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/XI0/N3
+ XI0/XI1/XI1/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=1.62e-13 AS=2.64e-13
+ PD=1.47e-06 PS=2.84e-06 M=1 sca=17.3113 scb=0.0168035 scc=0.00114318
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.03e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M4@4 XI0/XI1/XI1/N14 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/XI0/N3
+ XI0/XI1/XI1/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=1.62e-13 AS=2.64e-13
+ PD=1.47e-06 PS=2.84e-06 M=1 sca=7.68921 scb=0.0054437 scc=7.47049e-05
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.03e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M4@3 XI0/XI1/XI1/N14 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/XI0/N3
+ XI0/XI1/XI1/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=1.62e-13 AS=2.64e-13
+ PD=1.47e-06 PS=2.84e-06 M=1 sca=6.5521 scb=0.00532637 scc=7.46664e-05
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.03e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/XI0/M4@2 XI0/XI1/XI1/N14 XI0/XI1/XI1/XI0/N2 XI0/XI1/XI1/XI0/N3
+ XI0/XI1/XI1/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=1.62e-13 AS=2.64e-13
+ PD=1.47e-06 PS=2.84e-06 M=1 sca=9.16105 scb=0.00687439 scc=8.49142e-05
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.03e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M26 XI0/XI1/XI1/N9 XI0/XI1/XI1/N14 VSSA_TX VSSA_TX egnfet L=7e-07
+ W=4.6e-07 AD=6.21e-14 AS=1.012e-13 PD=7.3e-07 PS=1.36e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=2.2e-07 sb=1.19e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M26@2 XI0/XI1/XI1/N9 XI0/XI1/XI1/N14 VSSA_TX VSSA_TX egnfet L=7e-07
+ W=4.6e-07 AD=6.21e-14 AS=1.012e-13 PD=7.3e-07 PS=1.36e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=1.19e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M25 XI0/XI1/XI1/N10 XI0/XI1/XI1/N14 VSSA_TX VSSA_TX egnfet L=7e-07
+ W=4.6e-07 AD=6.21e-14 AS=1.012e-13 PD=7.3e-07 PS=1.36e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=2.2e-07 sb=1.19e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M25@2 XI0/XI1/XI1/N10 XI0/XI1/XI1/N14 VSSA_TX VSSA_TX egnfet
+ L=7e-07 W=4.6e-07 AD=6.21e-14 AS=1.012e-13 PD=7.3e-07 PS=1.36e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=1.19e-06 sb=2.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M18 XI0/XI1/XI1/N8 XI0/XI1/XI1/N8 XI0/XI1/XI1/N1N22 VSSA_TX egnfet
+ L=6e-07 W=6.2e-07 AD=1.364e-13 AS=8.37e-14 PD=1.68e-06 PS=8.9e-07 M=1
+ sca=0.960238 scb=4.29893e-05 scc=2.6802e-09 lpccnr=5.55e-07 covpccnr=0
+ wrxcnr=5.58e-07 sa=2.2e-07 sb=1.09e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M18@2 XI0/XI1/XI1/N8 XI0/XI1/XI1/N8 XI0/XI1/XI1/N1N22 VSSA_TX
+ egnfet L=6e-07 W=6.2e-07 AD=1.364e-13 AS=8.37e-14 PD=1.68e-06 PS=8.9e-07 M=1
+ sca=0.960238 scb=4.29893e-05 scc=2.6802e-09 lpccnr=5.55e-07 covpccnr=0
+ wrxcnr=5.58e-07 sa=1.09e-06 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M16 XI0/XI1/XI1/N1N22 XI0/XI1/XI1/N8 VSSA_TX VSSA_TX egnfet
+ L=1.2e-06 W=5e-07 AD=1.1e-13 AS=1.1e-13 PD=1.44e-06 PS=1.44e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=1.095e-06 covpccnr=0 wrxcnr=4.5e-07 sa=2.2e-07 sb=2.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M15 XI0/XI1/XI1/N1N24 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=2.2e-07 sb=1.09e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M17 XI0/XI1/XI1/N7 XI0/XI1/XI1/N8 XI0/XI1/XI1/N1N24 VSSA_TX egnfet
+ L=6e-07 W=1.54e-06 AD=3.388e-13 AS=2.079e-13 PD=3.52e-06 PS=1.81e-06 M=1
+ sca=0.72776 scb=1.92596e-05 scc=1.08865e-09 lpccnr=5.55e-07 covpccnr=0
+ wrxcnr=1.386e-06 sa=2.2e-07 sb=1.09e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M15@2 XI0/XI1/XI1/N1N24 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet
+ L=6e-07 W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=1.09e-06 sb=2.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M17@2 XI0/XI1/XI1/N7 XI0/XI1/XI1/N8 XI0/XI1/XI1/N1N24 VSSA_TX
+ egnfet L=6e-07 W=1.54e-06 AD=3.388e-13 AS=2.079e-13 PD=3.52e-06 PS=1.81e-06
+ M=1 sca=0.72776 scb=1.92596e-05 scc=1.08865e-09 lpccnr=5.55e-07 covpccnr=0
+ wrxcnr=1.386e-06 sa=1.09e-06 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M24 XI0/XI1/XI1/N9 XI0/XI1/XI1/N9 XI0/XI1/XI1/N1N21 VDDHA_TX egpfet
+ L=3e-07 W=1.88e-06 AD=4.136e-13 AS=2.538e-13 PD=4.2e-06 PS=2.15e-06 M=1
+ sca=7.74306 scb=0.00682578 scc=0.0001436 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=1.692e-06 sa=2.2e-07 sb=7.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M24@2 XI0/XI1/XI1/N9 XI0/XI1/XI1/N9 XI0/XI1/XI1/N1N21 VDDHA_TX
+ egpfet L=3e-07 W=1.88e-06 AD=4.136e-13 AS=2.538e-13 PD=4.2e-06 PS=2.15e-06 M=1
+ sca=5.71348 scb=0.00412582 scc=0.000121924 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=1.692e-06 sa=7.9e-07 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M22 XI0/XI1/XI1/N1N21 XI0/XI1/XI1/N9 VDDHA_TX VDDHA_TX egpfet
+ L=4e-07 W=7.2e-07 AD=1.584e-13 AS=1.584e-13 PD=1.88e-06 PS=1.88e-06 M=1
+ sca=1.7507 scb=0.000410856 scc=2.68924e-07 lpccnr=3.75e-07 covpccnr=0
+ wrxcnr=6.48e-07 sa=2.2e-07 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M23 XI0/XI1/XI1/N10 XI0/XI1/XI1/N9 XI0/XI1/XI1/N1N4 VDDHA_TX egpfet
+ L=3e-07 W=3.76e-06 AD=8.289e-13 AS=5.0845e-13 PD=7.98e-06 PS=4.04e-06 M=1
+ sca=2.21946 scb=0.00182982 scc=6.07933e-05 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.38401e-06 sa=2.2e-07 sb=7.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M23@2 XI0/XI1/XI1/N10 XI0/XI1/XI1/N9 XI0/XI1/XI1/N1N4 VDDHA_TX
+ egpfet L=3e-07 W=3.76e-06 AD=8.289e-13 AS=5.0845e-13 PD=7.98e-06 PS=4.04e-06
+ M=1 sca=2.21946 scb=0.00182982 scc=6.07933e-05 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.38401e-06 sa=7.9e-07 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M21 XI0/XI1/XI1/N1N4 XI0/XI1/XI1/N10 VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1
+ sca=1.89484 scb=0.000866238 scc=4.73755e-06 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=1.692e-06 sa=2.2e-07 sb=7.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M21@2 XI0/XI1/XI1/N1N4 XI0/XI1/XI1/N10 VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1
+ sca=1.89484 scb=0.000866238 scc=4.73755e-06 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=1.692e-06 sa=7.9e-07 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M19 XI0/XI1/XI1/N8 XI0/XI1/XI1/N10 VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1 sca=1.89484
+ scb=0.000866238 scc=4.73755e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06
+ sa=2.2e-07 sb=7.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M19@2 XI0/XI1/XI1/N8 XI0/XI1/XI1/N10 VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1
+ sca=1.89484 scb=0.000866238 scc=4.73755e-06 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=1.692e-06 sa=7.9e-07 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M20 XI0/XI1/XI1/N7 XI0/XI1/XI1/N10 VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1 sca=1.89484
+ scb=0.000866238 scc=4.73755e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06
+ sa=2.2e-07 sb=7.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M20@2 XI0/XI1/XI1/N7 XI0/XI1/XI1/N10 VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1
+ sca=1.89484 scb=0.000866238 scc=4.73755e-06 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=1.692e-06 sa=7.9e-07 sb=2.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M11 XI0/XI1/XI1/N1 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=2.2e-07 sb=1.09e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M11@6 XI0/XI1/XI1/N1 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=1.09e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M11@5 XI0/XI1/XI1/N1 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=2.2e-07 sb=1.09e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M11@4 XI0/XI1/XI1/N1 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=1.09e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M11@3 XI0/XI1/XI1/N1 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=2.2e-07 sb=1.09e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M11@2 XI0/XI1/XI1/N1 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=1.09e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M5@2 XI0/XI1/XI1/N4 XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.93e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/MD@3 VDDHA_TX VDDHA_TX VDDHA_TX VDDHA_TX egpfet L=2.8e-07 W=4e-06
+ AD=8.8e-13 AS=8.8e-13 PD=8.44e-06 PS=8.44e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.2e-07 sb=2.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M1@9 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet L=2.8e-07
+ W=4e-06 AD=5.4e-13 AS=8.8e-13 PD=4.27e-06 PS=8.44e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M1@8 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet L=2.8e-07
+ W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=7.7e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M1@7 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet L=2.8e-07
+ W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.32e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M1@6 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet L=2.8e-07
+ W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.87e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M1@5 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet L=2.8e-07
+ W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=1.87e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M1@4 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet L=2.8e-07
+ W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=1.32e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M3 XI0/XI1/XI1/N3 XI0/XI1/XI1/N10 VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=2.2e-07 sb=7.9e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M1@3 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet L=2.8e-07
+ W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=7.7e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M1@2 XI0/XI1/XI1/N1 XI0/FB XI0/XI1/XI1/N3 VDDHA_TX egpfet L=2.8e-07
+ W=4e-06 AD=5.4e-13 AS=8.8e-13 PD=4.27e-06 PS=8.44e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M3@4 XI0/XI1/XI1/N3 XI0/XI1/XI1/N10 VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=7.9e-07 sb=2.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M12 XI0/XI1/XI1/N2 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=2.2e-07 sb=1.09e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M12@6 XI0/XI1/XI1/N2 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=1.09e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M12@5 XI0/XI1/XI1/N2 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=2.2e-07 sb=1.09e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M12@4 XI0/XI1/XI1/N2 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=1.09e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M12@3 XI0/XI1/XI1/N2 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=2.2e-07 sb=1.09e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M12@2 XI0/XI1/XI1/N2 XI0/XI1/XI1/N7 VSSA_TX VSSA_TX egnfet L=6e-07
+ W=6.2e-07 AD=8.37e-14 AS=1.364e-13 PD=8.9e-07 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=1.09e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M6@2 XI0/XI1/XI1/N5 XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.93e-06 sb=2.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/MD@2 VDDHA_TX VDDHA_TX VDDHA_TX VDDHA_TX egpfet L=2.8e-07 W=4e-06
+ AD=8.8e-13 AS=8.8e-13 PD=8.44e-06 PS=8.44e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.2e-07 sb=2.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2@9 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=8.8e-13 PD=4.27e-06 PS=8.44e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.2e-07 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M2@8 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=7.7e-07 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M2@7 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.32e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2@6 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.87e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2@5 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06
+ sb=1.87e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M2@4 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06
+ sb=1.32e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M3@3 XI0/XI1/XI1/N3 XI0/XI1/XI1/N10 VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=2.2e-07 sb=7.9e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M2@3 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=5.4e-13 PD=4.27e-06 PS=4.27e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=7.7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M2@2 XI0/XI1/XI1/N2 XI0/VCM XI0/XI1/XI1/N3 VDDHA_TX egpfet
+ L=2.8e-07 W=4e-06 AD=5.4e-13 AS=8.8e-13 PD=4.27e-06 PS=8.44e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=2.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M3@2 XI0/XI1/XI1/N3 XI0/XI1/XI1/N10 VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=1.88e-06 AD=2.538e-13 AS=4.136e-13 PD=2.15e-06 PS=4.2e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=7.9e-07 sb=2.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XI1/M27 VDDHA_TX XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=5e-06
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=6.58827
+ scb=0.00517796 scc=0.000563345 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M27@4 VDDHA_TX XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=5e-06
+ W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M27@3 VDDHA_TX XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=5e-06
+ W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=4.7619
+ scb=0.00367879 scc=0.000507507 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XI1/M27@2 VDDHA_TX XI0/XI1/XI1/N6 VDDHA_TX VDDHA_TX egpfet L=5e-06
+ W=5e-06 AD=6e-13 AS=3.5e-13 PD=1.024e-05 PS=5.14e-06 M=1 sca=10.5907
+ scb=0.00823657 scc=0.000989795 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XG1/M2 XI0/XI1/PD XI0/XI1/PDB VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07
+ AD=6.4e-14 AS=6.8e-14 PD=1.12e-06 PS=1.14e-06 M=1 sca=1.03966 scb=5.69875e-05
+ scc=3.99185e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.6e-07 sb=1.7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XG0/M2 XI0/XI1/PDB XI0/PDH VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07
+ AD=6.8e-14 AS=6.8e-14 PD=1.14e-06 PS=1.14e-06 M=1 sca=1.03966 scb=5.69875e-05
+ scc=3.99185e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.7e-07 sb=1.7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M26 XI0/VBP XI0/XI1/PDB VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1e-05
+ AD=1.1e-12 AS=1.7e-12 PD=1.022e-05 PS=2.034e-05 M=1 sca=1.2885 scb=0.000736082
+ scc=2.29206e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-06 sa=1.7e-07 sb=5.4e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/M26@2 XI0/VBP XI0/XI1/PDB VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1e-05
+ AD=1.1e-12 AS=1.7e-12 PD=1.022e-05 PS=2.034e-05 M=1 sca=1.2885 scb=0.000736082
+ scc=2.29206e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-06 sa=5.4e-07 sb=1.7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI1/XG1/M1 XI0/XI1/PD XI0/XI1/PDB VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=1.4e-06 AD=2.38e-13 AS=2.38e-13 PD=3.14e-06 PS=3.14e-06 M=1 sca=6.9286
+ scb=0.00560735 scc=0.000164091 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.7e-07 sb=1.7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI1/XG0/M1 XI0/XI1/PDB XI0/PDH VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=1.4e-06
+ AD=2.38e-13 AS=2.38e-13 PD=3.14e-06 PS=3.14e-06 M=1 sca=10.5958 scb=0.0114109
+ scc=0.000269279 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06 sa=1.7e-07
+ sb=1.7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XX287/X23/D0_noxref VSS VDD diodenwx  AREA=4.51385e-12 perim=8.85e-06 sizedup=0
XX287/X23/D1_noxref VSS VDD diodenwx  AREA=4.51385e-12 perim=8.85e-06 sizedup=0
XX287/X23/D2_noxref VSS VDD diodenwx  AREA=4.51385e-12 perim=8.85e-06 sizedup=0
XX287/X23/D3_noxref VSS VDD diodenwx  AREA=1.39566e-11 perim=1.553e-05 sizedup=0
XXI0/XI3A0/M4N XI0/XI3A0/N3 CCMI0 VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=1.08877 scb=6.77412e-05
+ scc=5.27538e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI3A1/M4N XI0/XI3A1/N3 CCMI1 VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=1.08877 scb=6.77412e-05
+ scc=5.27538e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI3A2/M4N XI0/XI3A2/N3 CCMI2 VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=1.08877 scb=6.77412e-05
+ scc=5.27538e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XG1/M2 XI0/N1N229 PDTXI VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=1.09334 scb=6.89641e-05
+ scc=5.47899e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XG2/M2 XI0/N1N225 XI0/N1N229 VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=1.09334 scb=6.89641e-05
+ scc=5.47899e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI2/M4N XI0/XI2/N3 XI0/N1N225 VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=1.08877 scb=6.77412e-05
+ scc=5.27538e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XG3/M2 XI0/EN XI0/N1N225 VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=1.09334 scb=6.89641e-05
+ scc=5.47899e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI3A0/XG2/M2 XI0/CCMH0 XI0/XI3A0/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/XG2/M2@4 XI0/CCMH0 XI0/XI3A0/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/XG2/M2@3 XI0/CCMH0 XI0/XI3A0/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/XG2/M2@2 XI0/CCMH0 XI0/XI3A0/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/XG1/M2 XI0/XI3A0/N1N36 XI0/XI3A0/N1N5 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06 M=1
+ sca=0.985416 scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=7.2e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/M4P XI0/XI3A0/N1N5 XI0/XI3A0/N2 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999
+ scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/M2P XI0/XI3A0/N2 CCMI0 VSSA_TX VSSA_TX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=1.04193
+ scb=6.22794e-05 scc=5.97817e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/M2N XI0/XI3A0/N1 XI0/XI3A0/N3 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=6.4e-07 AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=1.04193
+ scb=6.22794e-05 scc=5.97817e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/XG2/M2 XI0/CCMH1 XI0/XI3A1/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/XG2/M2@4 XI0/CCMH1 XI0/XI3A1/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/XG2/M2@3 XI0/CCMH1 XI0/XI3A1/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/XG2/M2@2 XI0/CCMH1 XI0/XI3A1/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/XG1/M2 XI0/XI3A1/N1N36 XI0/XI3A1/N1N5 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06 M=1
+ sca=0.985416 scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=7.2e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/M4P XI0/XI3A1/N1N5 XI0/XI3A1/N2 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999
+ scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/M2P XI0/XI3A1/N2 CCMI1 VSSA_TX VSSA_TX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=1.04193
+ scb=6.22794e-05 scc=5.97817e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/M2N XI0/XI3A1/N1 XI0/XI3A1/N3 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=6.4e-07 AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=1.04193
+ scb=6.22794e-05 scc=5.97817e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/XG2/M2 XI0/CCMH2 XI0/XI3A2/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/XG2/M2@4 XI0/CCMH2 XI0/XI3A2/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/XG2/M2@3 XI0/CCMH2 XI0/XI3A2/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/XG2/M2@2 XI0/CCMH2 XI0/XI3A2/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/XG1/M2 XI0/XI3A2/N1N36 XI0/XI3A2/N1N5 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06 M=1
+ sca=0.985416 scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=7.2e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/M4P XI0/XI3A2/N1N5 XI0/XI3A2/N2 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999
+ scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/M2P XI0/XI3A2/N2 CCMI2 VSSA_TX VSSA_TX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=1.04193
+ scb=6.22794e-05 scc=5.97817e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/M2N XI0/XI3A2/N1 XI0/XI3A2/N3 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=6.4e-07 AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=1.04193
+ scb=6.22794e-05 scc=5.97817e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI2/XG2/M2 XI0/PDH XI0/XI2/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0.985416 scb=5.22299e-05
+ scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=9.9e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI2/XG2/M2@4 XI0/PDH XI0/XI2/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0.985416 scb=5.22299e-05
+ scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI2/XG2/M2@3 XI0/PDH XI0/XI2/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0.985416 scb=5.22299e-05
+ scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=7e-07 sb=4.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI2/XG2/M2@2 XI0/PDH XI0/XI2/N1N36 VSSA_TX VSSA_TX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0.985416 scb=5.22299e-05
+ scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=9.9e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI2/XG1/M2 XI0/XI2/N1N36 XI0/XI2/N1N5 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06 M=1 sca=0.985416
+ scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI2/M4P XI0/XI2/N1N5 XI0/XI2/N2 VSSA_TX VSSA_TX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=1.13999 scb=8.44443e-05
+ scc=9.17689e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI2/M2P XI0/XI2/N2 XI0/N1N225 VSSA_TX VSSA_TX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=1.04193
+ scb=6.22794e-05 scc=5.97817e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI2/M2N XI0/XI2/N1 XI0/XI2/N3 VSSA_TX VSSA_TX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=1.04193
+ scb=6.22794e-05 scc=5.97817e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/M3N XI0/XI3A0/N3 CCMI0 VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=29.0869 scb=0.0336188
+ scc=0.00177331 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI3A1/M3N XI0/XI3A1/N3 CCMI1 VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=29.0869 scb=0.0336188
+ scc=0.00177331 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI3A2/M3N XI0/XI3A2/N3 CCMI2 VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=29.0869 scb=0.0336188
+ scc=0.00177331 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XG1/M1 XI0/N1N229 PDTXI VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=12.081 scb=0.0113715
+ scc=0.000401439 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XG2/M1 XI0/N1N225 XI0/N1N229 VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=11.4343 scb=0.0108379
+ scc=0.000400581 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI2/M3N XI0/XI2/N3 XI0/N1N225 VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=9.01787 scb=0.00609704
+ scc=5.7811e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XG3/M1 XI0/EN XI0/N1N225 VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=22.8249 scb=0.0278237
+ scc=0.0014721 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI3A0/XG2/M1 XI0/CCMH0 XI0/XI3A0/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=6.12186
+ scb=0.00459451 scc=0.000151456 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/XG2/M1@4 XI0/CCMH0 XI0/XI3A0/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=5.31379
+ scb=0.00369972 scc=0.000148393 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/XG2/M1@3 XI0/CCMH0 XI0/XI3A0/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=4.81796
+ scb=0.00336006 scc=0.000148032 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/XG2/M1@2 XI0/CCMH0 XI0/XI3A0/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=4.49198
+ scb=0.00323503 scc=0.000147991 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/XG1/M1 XI0/XI3A0/N1N36 XI0/XI3A0/N1N5 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=2.8e-06 AD=3.36e-13 AS=3.36e-13 PD=5.84e-06 PS=5.84e-06 M=1
+ sca=3.39213 scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.52e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/M3P XI0/XI3A0/N1N5 XI0/XI3A0/N2 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=3.32164
+ scb=0.00268154 scc=4.15811e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/M1P XI0/XI3A0/N2 XI0/XI3A0/N1 VDDHA_TX VDDHA_TX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.15302
+ scb=0.00156258 scc=3.15078e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A0/M1N XI0/XI3A0/N1 XI0/XI3A0/N2 VDDHA_TX VDDHA_TX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.15302
+ scb=0.00156258 scc=3.15078e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/XG2/M1 XI0/CCMH1 XI0/XI3A1/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/XG2/M1@4 XI0/CCMH1 XI0/XI3A1/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/XG2/M1@3 XI0/CCMH1 XI0/XI3A1/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/XG2/M1@2 XI0/CCMH1 XI0/XI3A1/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/XG1/M1 XI0/XI3A1/N1N36 XI0/XI3A1/N1N5 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=2.8e-06 AD=3.36e-13 AS=3.36e-13 PD=5.84e-06 PS=5.84e-06 M=1
+ sca=3.39213 scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.52e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/M3P XI0/XI3A1/N1N5 XI0/XI3A1/N2 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=3.32164
+ scb=0.00268154 scc=4.15811e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/M1P XI0/XI3A1/N2 XI0/XI3A1/N1 VDDHA_TX VDDHA_TX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.15302
+ scb=0.00156258 scc=3.15078e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A1/M1N XI0/XI3A1/N1 XI0/XI3A1/N2 VDDHA_TX VDDHA_TX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.15302
+ scb=0.00156258 scc=3.15078e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/XG2/M1 XI0/CCMH2 XI0/XI3A2/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/XG2/M1@4 XI0/CCMH2 XI0/XI3A2/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/XG2/M1@3 XI0/CCMH2 XI0/XI3A2/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/XG2/M1@2 XI0/CCMH2 XI0/XI3A2/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/XG1/M1 XI0/XI3A2/N1N36 XI0/XI3A2/N1N5 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=2.8e-06 AD=3.36e-13 AS=3.36e-13 PD=5.84e-06 PS=5.84e-06 M=1
+ sca=3.39213 scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.52e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/M3P XI0/XI3A2/N1N5 XI0/XI3A2/N2 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=3.32164
+ scb=0.00268154 scc=4.15811e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/M1P XI0/XI3A2/N2 XI0/XI3A2/N1 VDDHA_TX VDDHA_TX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.15302
+ scb=0.00156258 scc=3.15078e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI3A2/M1N XI0/XI3A2/N1 XI0/XI3A2/N2 VDDHA_TX VDDHA_TX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.15302
+ scb=0.00156258 scc=3.15078e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI2/XG2/M1 XI0/PDH XI0/XI2/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI2/XG2/M1@4 XI0/PDH XI0/XI2/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI2/XG2/M1@3 XI0/PDH XI0/XI2/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI2/XG2/M1@2 XI0/PDH XI0/XI2/N1N36 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI2/XG1/M1 XI0/XI2/N1N36 XI0/XI2/N1N5 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=2.8e-06 AD=3.36e-13 AS=3.36e-13 PD=5.84e-06 PS=5.84e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI2/M3P XI0/XI2/N1N5 XI0/XI2/N2 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=3.32164
+ scb=0.00268154 scc=4.15811e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI2/M1P XI0/XI2/N2 XI0/XI2/N1 VDDHA_TX VDDHA_TX egpfet L=3e-06 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.15302 scb=0.00156258
+ scc=3.15078e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI2/M1N XI0/XI2/N1 XI0/XI2/N2 VDDHA_TX VDDHA_TX egpfet L=3e-06 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=4.25724 scb=0.00228655
+ scc=3.24226e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XX287/X24/D0_noxref VSS VDD diodenwx  AREA=4.51385e-12 perim=8.85e-06 sizedup=0
XX287/X24/D1_noxref VSS VDDHA_TX diodenwx  AREA=1.53962e-10 perim=5.79e-05
+ sizedup=0
XX287/X24/D2_noxref VSS VDDHA_TX diodenwx  AREA=3.48534e-10 perim=0.00010642
+ sizedup=0
XX287/X24/D3_noxref VSS VDDHA_TX diodenwx  AREA=2.52916e-09 perim=0.00031288
+ sizedup=0
XXI0/XI0/XI2/X1I43/M4N XI0/XI0/XI2/X1I43/N3 XI0/EN VSS VSS nfet L=3e-08
+ W=2.8e-07 AD=2.94e-14 AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=1.08877
+ scb=6.77412e-05 scc=5.27538e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/M2N XI0/XI0/XI2/X1I43/N1 XI0/XI0/XI2/X1I43/N3 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=6.4e-07 AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1
+ sca=1.04193 scb=6.22794e-05 scc=5.97817e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/M2P XI0/XI0/XI2/X1I43/N2 XI0/EN VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=6.4e-07 AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1
+ sca=1.04193 scb=6.22794e-05 scc=5.97817e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/M4P XI0/XI0/XI2/X1I43/N1N5 XI0/XI0/XI2/X1I43/N2 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06
+ M=1 sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/XG1/M2 XI0/XI0/XI2/X1I43/N1N36 XI0/XI0/XI2/X1I43/N1N5 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06
+ M=1 sca=0.985416 scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=7.2e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/XG2/M2 XI0/XI0/XI2/PDB XI0/XI0/XI2/X1I43/N1N36 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06
+ M=1 sca=0.985416 scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=7.2e-07 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/XG2/M2@4 XI0/XI0/XI2/PDB XI0/XI0/XI2/X1I43/N1N36 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07
+ M=1 sca=0.985416 scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=7.2e-07 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/XG2/M2@3 XI0/XI0/XI2/PDB XI0/XI0/XI2/X1I43/N1N36 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07
+ M=1 sca=0.985416 scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=7.2e-07 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/XG2/M2@2 XI0/XI0/XI2/PDB XI0/XI0/XI2/X1I43/N1N36 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06
+ M=1 sca=0.985416 scb=5.22299e-05 scc=4.80861e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=7.2e-07 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/M3N XI0/XI0/XI2/X1I43/N3 XI0/EN VDD VDD pfet L=3e-08
+ W=5.6e-07 AD=5.88e-14 AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=29.0869
+ scb=0.0336188 scc=0.00177331 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/M1N XI0/XI0/XI2/X1I43/N1 XI0/XI0/XI2/X1I43/N2 VDDHA_TX
+ VDDHA_TX egpfet L=3e-06 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06
+ M=1 sca=4.25724 scb=0.00228655 scc=3.24226e-05 lpccnr=2.715e-06 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/M1P XI0/XI0/XI2/X1I43/N2 XI0/XI0/XI2/X1I43/N1 VDDHA_TX
+ VDDHA_TX egpfet L=3e-06 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06
+ M=1 sca=2.15302 scb=0.00156258 scc=3.15078e-05 lpccnr=2.715e-06 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/M3P XI0/XI0/XI2/X1I43/N1N5 XI0/XI0/XI2/X1I43/N2 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06
+ PS=3.04e-06 M=1 sca=3.32164 scb=0.00268154 scc=4.15811e-05 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/XG1/M1 XI0/XI0/XI2/X1I43/N1N36 XI0/XI0/XI2/X1I43/N1N5
+ VDDHA_TX VDDHA_TX egpfet L=1.5e-07 W=2.8e-06 AD=3.36e-13 AS=3.36e-13
+ PD=5.84e-06 PS=5.84e-06 M=1 sca=3.39213 scb=0.00316561 scc=0.000147986
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/XG2/M1 XI0/XI0/XI2/PDB XI0/XI0/XI2/X1I43/N1N36 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06
+ PS=5.84e-06 M=1 sca=3.39213 scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=2.52e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/XG2/M1@4 XI0/XI0/XI2/PDB XI0/XI0/XI2/X1I43/N1N36 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06
+ PS=2.94e-06 M=1 sca=3.39213 scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=2.52e-06 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/XG2/M1@3 XI0/XI0/XI2/PDB XI0/XI0/XI2/X1I43/N1N36 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06
+ PS=2.94e-06 M=1 sca=3.39213 scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=2.52e-06 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I43/XG2/M1@2 XI0/XI0/XI2/PDB XI0/XI0/XI2/X1I43/N1N36 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06
+ PS=5.84e-06 M=1 sca=3.39213 scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=2.52e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XX287/X24/X24/D0_noxref VSS VDD diodenwx  AREA=7.95448e-11 perim=4.724e-05
+ sizedup=0
XXI0/XI0/XI3/X1I221/M0 XI0/XI0/XI3/X1I221/N1N42 XI0/XI0/XI3/X1I221/N1N42 VSS VSS
+ nfet L=3e-08 W=1.1e-07 AD=2.09e-14 AS=2.09e-14 PD=6e-07 PS=6e-07 M=1
+ sca=1.77931 scb=0.000417271 scc=2.35895e-07 lpccnr=3.1e-08 covpccnr=0
+ wrxcnr=9.9e-08 sa=1.9e-07 sb=1.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG12/M2 XI0/XI0/NP1 XI0/XI0/XI3/N1N206 VSS VSS nfet L=3e-08 W=7e-07
+ AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=1.36272 scb=0.000187218
+ scc=6.5656e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07 sa=1.05e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG12/M2@4 XI0/XI0/NP1 XI0/XI0/XI3/N1N206 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=1.36272
+ scb=0.000187218 scc=6.5656e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=2.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG12/M2@3 XI0/XI0/NP1 XI0/XI0/XI3/N1N206 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=1.36272
+ scb=0.000187218 scc=6.5656e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=4.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG12/M2@2 XI0/XI0/NP1 XI0/XI0/XI3/N1N206 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=1.36272
+ scb=0.000187218 scc=6.5656e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=5.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG11/M4 XI0/XI0/XI3/XG11/N1 XI0/EN VSS VSS nfet L=3e-08 W=1.4e-06
+ AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=1.06648 scb=0.000101269
+ scc=3.29931e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06 sa=1.05e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG11/M3 XI0/XI0/XI3/N1N206 XI0/XI0/XI3/N0P XI0/XI0/XI3/XG11/N1 VSS
+ nfet L=3e-08 W=1.4e-06 AD=1.47e-13 AS=8.4e-14 PD=3.01e-06 PS=1.52e-06 M=1
+ sca=1.06648 scb=0.000101269 scc=3.29931e-08 lpccnr=3.1e-08 covpccnr=0
+ wrxcnr=1.26e-06 sa=2.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG6/M2 XI0/XI0/XI3/N0P XI0/XI0/XI3/NN VSS VSS nfet L=3e-08
+ W=3.5e-07 AD=2.1e-14 AS=3.675e-14 PD=4.7e-07 PS=9.1e-07 M=1 sca=1.58252
+ scb=0.000290095 scc=1.22506e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.15e-07
+ sa=1.05e-07 sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG6/M2@4 XI0/XI0/XI3/N0P XI0/XI0/XI3/NN VSS VSS nfet L=3e-08
+ W=3.5e-07 AD=2.1e-14 AS=2.1e-14 PD=4.7e-07 PS=4.7e-07 M=1 sca=1.58252
+ scb=0.000290095 scc=1.22506e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.15e-07
+ sa=2.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG6/M2@3 XI0/XI0/XI3/N0P XI0/XI0/XI3/NN VSS VSS nfet L=3e-08
+ W=3.5e-07 AD=2.1e-14 AS=2.1e-14 PD=4.7e-07 PS=4.7e-07 M=1 sca=1.58252
+ scb=0.000290095 scc=1.22506e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.15e-07
+ sa=4.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG6/M2@2 XI0/XI0/XI3/N0P XI0/XI0/XI3/NN VSS VSS nfet L=3e-08
+ W=3.5e-07 AD=2.1e-14 AS=3.675e-14 PD=4.7e-07 PS=9.1e-07 M=1 sca=1.58252
+ scb=0.000290095 scc=1.22506e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.15e-07
+ sa=5.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG7/M2 XI0/XI0/XI3/N0N XI0/XI0/XI3/NP VSS VSS nfet L=3e-08
+ W=3.5e-07 AD=2.1e-14 AS=3.675e-14 PD=4.7e-07 PS=9.1e-07 M=1 sca=1.58252
+ scb=0.000290095 scc=1.22506e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.15e-07
+ sa=1.05e-07 sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG7/M2@4 XI0/XI0/XI3/N0N XI0/XI0/XI3/NP VSS VSS nfet L=3e-08
+ W=3.5e-07 AD=2.1e-14 AS=2.1e-14 PD=4.7e-07 PS=4.7e-07 M=1 sca=1.58252
+ scb=0.000290095 scc=1.22506e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.15e-07
+ sa=2.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG7/M2@3 XI0/XI0/XI3/N0N XI0/XI0/XI3/NP VSS VSS nfet L=3e-08
+ W=3.5e-07 AD=2.1e-14 AS=2.1e-14 PD=4.7e-07 PS=4.7e-07 M=1 sca=1.58252
+ scb=0.000290095 scc=1.22506e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.15e-07
+ sa=4.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG7/M2@2 XI0/XI0/XI3/N0N XI0/XI0/XI3/NP VSS VSS nfet L=3e-08
+ W=3.5e-07 AD=2.1e-14 AS=3.675e-14 PD=4.7e-07 PS=9.1e-07 M=1 sca=1.58252
+ scb=0.000290095 scc=1.22506e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.15e-07
+ sa=5.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG10/M3 XI0/XI0/XI3/N1N207 XI0/XI0/XI3/N0N XI0/XI0/XI3/XG10/N1 VSS
+ nfet L=3e-08 W=1.4e-06 AD=1.47e-13 AS=8.4e-14 PD=3.01e-06 PS=1.52e-06 M=1
+ sca=1.06648 scb=0.000101269 scc=3.29931e-08 lpccnr=3.1e-08 covpccnr=0
+ wrxcnr=1.26e-06 sa=1.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG10/M4 XI0/XI0/XI3/XG10/N1 XI0/EN VSS VSS nfet L=3e-08 W=1.4e-06
+ AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=1.06648 scb=0.000101269
+ scc=3.29931e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06 sa=2.55e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG13/M2 XI0/XI0/NN1 XI0/XI0/XI3/N1N207 VSS VSS nfet L=3e-08 W=7e-07
+ AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=2.39976 scb=0.000240619
+ scc=6.85634e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07 sa=1.05e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG13/M2@4 XI0/XI0/NN1 XI0/XI0/XI3/N1N207 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=2.53913
+ scb=0.000278574 scc=7.4719e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=2.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG13/M2@3 XI0/XI0/NN1 XI0/XI0/XI3/N1N207 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=2.70861
+ scb=0.000342846 scc=9.37874e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=4.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG13/M2@2 XI0/XI0/NN1 XI0/XI0/XI3/N1N207 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=2.91753
+ scb=0.00045105 scc=1.52553e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=5.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/X1I218/M0 XI0/XI0/XI3/TIEL XI0/XI0/XI3/X1I218/N1N50 VSS VSS nfet
+ L=3e-08 W=1.1e-07 AD=2.09e-14 AS=2.09e-14 PD=6e-07 PS=6e-07 M=1 sca=6.23088
+ scb=0.00456083 scc=3.6501e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9.9e-08
+ sa=1.9e-07 sb=1.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/X1I221/M1 XI0/XI0/XI3/TIEH XI0/XI0/XI3/X1I221/N1N42 VDD VDD pfet
+ L=3e-08 W=1.1e-07 AD=2.09e-14 AS=2.09e-14 PD=6e-07 PS=6e-07 M=1 sca=17.9968
+ scb=0.022339 scc=0.00116034 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9.9e-08
+ sa=1.9e-07 sb=1.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG12/M1 XI0/XI0/NP1 XI0/XI0/XI3/N1N206 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=5.63509
+ scb=0.0022769 scc=9.0426e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.05e-07 sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG12/M1@4 XI0/XI0/NP1 XI0/XI0/XI3/N1N206 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=5.25527
+ scb=0.00189176 scc=8.09045e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=2.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG12/M1@3 XI0/XI0/NP1 XI0/XI0/XI3/N1N206 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=4.96052
+ scb=0.00165848 scc=7.77618e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=4.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG12/M1@2 XI0/XI0/NP1 XI0/XI0/XI3/N1N206 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=4.72722
+ scb=0.00151843 scc=7.67324e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=5.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG11/M2 XI0/XI0/XI3/N1N206 XI0/EN VDD VDD pfet L=3e-08 W=1.4e-06
+ AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=3.28252 scb=0.00131567
+ scc=7.62377e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06 sa=1.05e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG11/M1 XI0/XI0/XI3/N1N206 XI0/XI0/XI3/N0P VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=3.28252
+ scb=0.00131567 scc=7.62377e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=2.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG6/M1 XI0/XI0/XI3/N0P XI0/XI0/XI3/NN VDD VDD pfet L=3e-08 W=7e-07
+ AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=3.25114 scb=0.00229244
+ scc=1.51359e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07 sa=1.05e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG6/M1@4 XI0/XI0/XI3/N0P XI0/XI0/XI3/NN VDD VDD pfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=3.25114
+ scb=0.00229244 scc=1.51359e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=2.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG6/M1@3 XI0/XI0/XI3/N0P XI0/XI0/XI3/NN VDD VDD pfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=3.25114
+ scb=0.00229244 scc=1.51359e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=4.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG8/M1 XI0/XI0/XI3/N0N XI0/XI0/XI3/N0P VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=1.47e-13 AS=1.47e-13 PD=3.01e-06 PS=3.01e-06 M=1 sca=4.68113
+ scb=0.00364992 scc=8.29514e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG6/M1@2 XI0/XI0/XI3/N0P XI0/XI0/XI3/NN VDD VDD pfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=3.25114
+ scb=0.00229244 scc=1.51359e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=5.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG7/M1 XI0/XI0/XI3/N0N XI0/XI0/XI3/NP VDD VDD pfet L=3e-08 W=7e-07
+ AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=3.25114 scb=0.00229244
+ scc=1.51359e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07 sa=1.05e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG9/M1 XI0/XI0/XI3/N0P XI0/XI0/XI3/N0N VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=1.47e-13 AS=1.47e-13 PD=3.01e-06 PS=3.01e-06 M=1 sca=4.68113
+ scb=0.00364992 scc=8.29514e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG7/M1@4 XI0/XI0/XI3/N0N XI0/XI0/XI3/NP VDD VDD pfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=3.25114
+ scb=0.00229244 scc=1.51359e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=2.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG7/M1@3 XI0/XI0/XI3/N0N XI0/XI0/XI3/NP VDD VDD pfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=3.25114
+ scb=0.00229244 scc=1.51359e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=4.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG7/M1@2 XI0/XI0/XI3/N0N XI0/XI0/XI3/NP VDD VDD pfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=3.25114
+ scb=0.00229244 scc=1.51359e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=5.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG10/M1 XI0/XI0/XI3/N1N207 XI0/XI0/XI3/N0N VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=3.28252
+ scb=0.00131567 scc=7.62377e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG10/M2 XI0/XI0/XI3/N1N207 XI0/EN VDD VDD pfet L=3e-08 W=1.4e-06
+ AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=3.28252 scb=0.00131567
+ scc=7.62377e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06 sa=2.55e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG13/M1 XI0/XI0/NN1 XI0/XI0/XI3/N1N207 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=4.72722
+ scb=0.00151843 scc=7.67324e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.05e-07 sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG13/M1@4 XI0/XI0/NN1 XI0/XI0/XI3/N1N207 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=4.96052
+ scb=0.00165848 scc=7.77618e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=2.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG13/M1@3 XI0/XI0/NN1 XI0/XI0/XI3/N1N207 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=5.25527
+ scb=0.00189176 scc=8.09045e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=4.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG13/M1@2 XI0/XI0/NN1 XI0/XI0/XI3/N1N207 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=5.63509
+ scb=0.0022769 scc=9.0426e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=5.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/X1I218/M1 XI0/XI0/XI3/X1I218/N1N50 XI0/XI0/XI3/X1I218/N1N50 VDD VDD
+ pfet L=3e-08 W=1.1e-07 AD=2.09e-14 AS=2.09e-14 PD=6e-07 PS=6e-07 M=1
+ sca=14.3923 scb=0.0175596 scc=0.00055081 lpccnr=3.1e-08 covpccnr=0
+ wrxcnr=9.9e-08 sa=1.9e-07 sb=1.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG8/M2 XI0/XI0/XI3/N0N XI0/XI0/XI3/N0P VSS VSS nfet L=3e-08 W=7e-07
+ AD=7.35e-14 AS=7.35e-14 PD=1.61e-06 PS=1.61e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG9/M2 XI0/XI0/XI3/N0P XI0/XI0/XI3/N0N VSS VSS nfet L=3e-08 W=7e-07
+ AD=7.35e-14 AS=7.35e-14 PD=1.61e-06 PS=1.61e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/MN XI0/XI0/XI3/IN4 XI0/XI0/XI3/TIEH XI0/XI0/XI3/NP VSS nfet L=3e-08
+ W=7e-07 AD=7.35e-14 AS=7.35e-14 PD=1.61e-06 PS=1.61e-06 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG1/M3 XI0/XI0/XI3/IN1 DTX XI0/XI0/XI3/XG1/N1 VSS nfet L=3e-08
+ W=4e-07 AD=4.2e-14 AS=2.4e-14 PD=1.01e-06 PS=5.2e-07 M=1 sca=1.03966
+ scb=5.69875e-05 scc=3.99185e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG1/M4 XI0/XI0/XI3/XG1/N1 XI0/EN VSS VSS nfet L=3e-08 W=4e-07
+ AD=2.4e-14 AS=4.2e-14 PD=5.2e-07 PS=1.01e-06 M=1 sca=1.03966 scb=5.69875e-05
+ scc=3.99185e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.6e-07 sa=2.55e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG2/M2 XI0/XI0/XI3/IN2 XI0/XI0/XI3/IN1 VSS VSS nfet L=3e-08 W=7e-07
+ AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=0.934286 scb=3.92097e-05
+ scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07 sa=1.05e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG2/M2@2 XI0/XI0/XI3/IN2 XI0/XI0/XI3/IN1 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=2.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG3/M2 XI0/XI0/XI3/IN3 XI0/XI0/XI3/IN2 VSS VSS nfet L=3e-08 W=7e-07
+ AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=0.934286 scb=3.92097e-05
+ scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07 sa=1.05e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG3/M2@4 XI0/XI0/XI3/IN3 XI0/XI0/XI3/IN2 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=2.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG3/M2@3 XI0/XI0/XI3/IN3 XI0/XI0/XI3/IN2 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=4.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG3/M2@2 XI0/XI0/XI3/IN3 XI0/XI0/XI3/IN2 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=5.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M2 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VSS VSS nfet L=3e-08 W=7e-07
+ AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=0.934286 scb=3.92097e-05
+ scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07 sa=1.05e-07
+ sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M2@8 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=2.55e-07 sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M2@7 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=4.05e-07 sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M2@6 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=5.55e-07 sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M2@5 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=7.05e-07 sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M2@4 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=8.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M2@3 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=1.005e-06 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M2@2 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=1.155e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG5/M2 XI0/XI0/XI3/NN XI0/XI0/XI3/IN4 VSS VSS nfet L=3e-08 W=7e-07
+ AD=4.2e-14 AS=7.35e-14 PD=8.2e-07 PS=1.61e-06 M=1 sca=0.934286 scb=3.92097e-05
+ scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07 sa=1.05e-07
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG5/M2@3 XI0/XI0/XI3/NN XI0/XI0/XI3/IN4 VSS VSS nfet L=3e-08
+ W=7e-07 AD=4.2e-14 AS=4.2e-14 PD=8.2e-07 PS=8.2e-07 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=2.55e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG5/M2@2 XI0/XI0/XI3/NN XI0/XI0/XI3/IN4 VSS VSS nfet L=3e-08
+ W=7e-07 AD=7.35e-14 AS=4.2e-14 PD=1.61e-06 PS=8.2e-07 M=1 sca=0.934286
+ scb=3.92097e-05 scc=2.3836e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=6.3e-07
+ sa=4.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/MP XI0/XI0/XI3/IN4 XI0/XI0/XI3/TIEL XI0/XI0/XI3/NP VDD pfet L=3e-08
+ W=1.4e-06 AD=1.47e-13 AS=1.47e-13 PD=3.01e-06 PS=3.01e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG1/M1 XI0/XI0/XI3/IN1 DTX VDD VDD pfet L=3e-08 W=4e-07 AD=2.4e-14
+ AS=4.2e-14 PD=5.2e-07 PS=1.01e-06 M=1 sca=9.39002 scb=0.0121669
+ scc=0.000535984 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.6e-07 sa=1.05e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG1/M2 XI0/XI0/XI3/IN1 XI0/EN VDD VDD pfet L=3e-08 W=4e-07
+ AD=2.4e-14 AS=4.2e-14 PD=5.2e-07 PS=1.01e-06 M=1 sca=9.39002 scb=0.0121669
+ scc=0.000535984 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.6e-07 sa=2.55e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG2/M1 XI0/XI0/XI3/IN2 XI0/XI0/XI3/IN1 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG2/M1@2 XI0/XI0/XI3/IN2 XI0/XI0/XI3/IN1 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=2.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG3/M1 XI0/XI0/XI3/IN3 XI0/XI0/XI3/IN2 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.05e-07 sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG3/M1@4 XI0/XI0/XI3/IN3 XI0/XI0/XI3/IN2 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=2.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG3/M1@3 XI0/XI0/XI3/IN3 XI0/XI0/XI3/IN2 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=4.05e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG3/M1@2 XI0/XI0/XI3/IN3 XI0/XI0/XI3/IN2 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=5.55e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M1 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.05e-07 sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M1@8 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=2.55e-07 sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M1@7 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=4.05e-07 sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M1@6 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=5.55e-07 sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M1@5 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=7.05e-07 sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M1@4 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=8.55e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M1@3 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.005e-06 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG4/M1@2 XI0/XI0/XI3/IN4 XI0/XI0/XI3/IN3 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.155e-06 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG5/M1 XI0/XI0/XI3/NN XI0/XI0/XI3/IN4 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=1.47e-13 PD=1.52e-06 PS=3.01e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.05e-07 sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG5/M1@3 XI0/XI0/XI3/NN XI0/XI0/XI3/IN4 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=8.4e-14 AS=8.4e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=2.55e-07 sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI3/XG5/M1@2 XI0/XI0/XI3/NN XI0/XI0/XI3/IN4 VDD VDD pfet L=3e-08
+ W=1.4e-06 AD=1.47e-13 AS=8.4e-14 PD=3.01e-06 PS=1.52e-06 M=1 sca=5.73611
+ scb=0.00492938 scc=0.000163279 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.26e-06
+ sa=4.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I45/M2 XI0/XI0/ENBH XI0/XI0/XI2/PDB VSSA_TX VSSA_TX egnfet
+ L=3.5e-07 W=8.4e-07 AD=1.008e-13 AS=1.008e-13 PD=1.92e-06 PS=1.92e-06 M=1
+ sca=0.972233 scb=5.0135e-05 scc=4.58236e-09 lpccnr=3.3e-07 covpccnr=0
+ wrxcnr=7.56e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M3 XI0/XI0/XI2/N1 XI0/XI0/NP1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1.25e-06 AD=8.75e-14 AS=1.5e-13 PD=1.39e-06 PS=2.74e-06 M=1 sca=1.85219
+ scb=0.000129326 scc=3.75783e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.125e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M3@2 XI0/XI0/XI2/N1 XI0/XI0/NP1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1.25e-06 AD=8.75e-14 AS=1.5e-13 PD=1.39e-06 PS=2.74e-06 M=1 sca=1.85219
+ scb=0.000129326 scc=3.75783e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.125e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M4 XI0/XI0/NP2 XI0/XI0/NN1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1.25e-06 AD=8.75e-14 AS=1.5e-13 PD=1.39e-06 PS=2.74e-06 M=1 sca=1.85219
+ scb=0.000129326 scc=3.75783e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.125e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M4@2 XI0/XI0/NP2 XI0/XI0/NN1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1.25e-06 AD=8.75e-14 AS=1.5e-13 PD=1.39e-06 PS=2.74e-06 M=1 sca=1.85219
+ scb=0.000129326 scc=3.75783e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.125e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M10 XI0/XI0/NN2 XI0/XI0/ENBH VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=1.23884
+ scb=0.000118379 scc=1.87971e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M8 XI0/XI0/NN2 XI0/XI0/NP1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1.25e-06 AD=8.75e-14 AS=1.5e-13 PD=1.39e-06 PS=2.74e-06 M=1 sca=1.85219
+ scb=0.000129326 scc=3.75783e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.125e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M8@2 XI0/XI0/NN2 XI0/XI0/NP1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1.25e-06 AD=8.75e-14 AS=1.5e-13 PD=1.39e-06 PS=2.74e-06 M=1 sca=1.85219
+ scb=0.000129326 scc=3.75783e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.125e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M7 XI0/XI0/XI2/N2 XI0/XI0/NN1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1.25e-06 AD=8.75e-14 AS=1.5e-13 PD=1.39e-06 PS=2.74e-06 M=1 sca=1.85219
+ scb=0.000129326 scc=3.75783e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.125e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M7@2 XI0/XI0/XI2/N2 XI0/XI0/NN1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1.25e-06 AD=8.75e-14 AS=1.5e-13 PD=1.39e-06 PS=2.74e-06 M=1 sca=1.85219
+ scb=0.000129326 scc=3.75783e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.125e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/X1I45/M1 XI0/XI0/ENBH XI0/XI0/XI2/PDB VDDHA_TX VDDHA_TX egpfet
+ L=3.5e-07 W=8.4e-07 AD=1.008e-13 AS=1.008e-13 PD=1.92e-06 PS=1.92e-06 M=1
+ sca=8.17528 scb=0.00980125 scc=0.00049195 lpccnr=3.3e-07 covpccnr=0
+ wrxcnr=7.56e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M11 XI0/XI0/XI2/N1 XI0/XI0/XI2/PDB VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=3.67129 scb=0.00286918 scc=1.89128e-05 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M1 XI0/XI0/XI2/N1 XI0/XI0/XI2/N1 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.98934
+ scb=0.000915443 scc=1.35474e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M1@2 XI0/XI0/XI2/N1 XI0/XI0/XI2/N1 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.98934
+ scb=0.000915443 scc=1.35474e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M2 XI0/XI0/NP2 XI0/XI0/XI2/N1 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.98934
+ scb=0.000915443 scc=1.35474e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M2@2 XI0/XI0/NP2 XI0/XI0/XI2/N1 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.98934
+ scb=0.000915443 scc=1.35474e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M9 XI0/XI0/NP2 XI0/XI0/XI2/PDB VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=3.67129
+ scb=0.00286918 scc=1.89128e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M6 XI0/XI0/NN2 XI0/XI0/XI2/N2 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.98934
+ scb=0.000915443 scc=1.35474e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M6@2 XI0/XI0/NN2 XI0/XI0/XI2/N2 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=1.98934
+ scb=0.000915443 scc=1.35474e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M5 XI0/XI0/XI2/N2 XI0/XI0/XI2/N2 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=3.17207
+ scb=0.00100949 scc=1.35573e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M5@2 XI0/XI0/XI2/N2 XI0/XI0/XI2/N2 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=3.53849
+ scb=0.00117751 scc=1.36354e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.5e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI2/M12 XI0/XI0/XI2/N2 XI0/XI0/XI2/PDB VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=9.36929 scb=0.00921682 scc=0.000117728 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XX287/X24/X35/D0_noxref VSS VDDHA_TX diodenwx  AREA=1.3844e-10 perim=5.645e-05
+ sizedup=0
XX287/X24/X35/D1_noxref VSS VDDHA_TX diodenwx  AREA=8.8008e-12 perim=1.228e-05
+ sizedup=0
XX287/X24/X35/D2_noxref VSS VDDHA_TX diodenwx  AREA=4.01512e-10 perim=0.00035532
+ sizedup=0
XX287/X24/X35/D3_noxref VSS XI0/XI0/XI0/XI0/N1 diodenwx  AREA=1.82161e-10
+ perim=6.394e-05 sizedup=0
XX287/X24/X35/D4_noxref VSS VDDHA_TX diodenwx  AREA=2.50573e-10 perim=8.238e-05
+ sizedup=0
XX287/X24/X35/D5_noxref VSS VDDHA_TX diodenwx  AREA=1.41514e-11 perim=1.51e-05
+ sizedup=0
XXI0/XI0/XI0/XI0/RRF XI0/XI0/CM XI0/XI0/XI0/XI0/N1N152 VDDHA_TX opppcres 231.017
+ M=1 w=2.945e-06 l=1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI0/XI0/RRC XI0/XI0/XI0/N3 XI0/XI0/XI0/VBN VDDHA_TX opppcres 968.268 M=1
+ w=2e-06 l=3.08e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI0/XI0/CC55 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC54 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC53 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC52 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC51 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC50 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC49 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC48 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC47 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC46 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC45 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC44 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC43 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC42 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC41 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC40 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC39 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC38 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC0 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC1 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC2 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC3 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC4 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC5 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC6 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC7 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC8 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC9 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC10 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC11 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC12 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC13 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC14 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC15 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC16 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC17 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC18 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC19 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC20 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC21 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC22 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC23 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC24 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC25 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC26 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC27 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC28 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC29 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC30 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC31 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC32 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC33 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC34 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC35 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC36 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/CC37 XI0/XI0/CM XI0/XI0/XI0/N3 VSSA_TX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI0/XI0/XI0/XI0/M9P XI0/XI0/XI0/XI0/N2N XI0/XI0/ENBH VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M3N XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N2N VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1
+ sca=1.66903 scb=0.000119808 scc=4.71809e-08 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M3N@2 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N2N VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1
+ sca=1.66903 scb=0.000119808 scc=4.71809e-08 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M3P XI0/XI0/XI0/VBN XI0/XI0/XI0/XI0/N2N VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1
+ sca=1.66903 scb=0.000119808 scc=4.71809e-08 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M3P@2 XI0/XI0/XI0/VBN XI0/XI0/XI0/XI0/N2N VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1
+ sca=1.66903 scb=0.000119808 scc=4.71809e-08 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M9N XI0/XI0/XI0/VBN XI0/XI0/ENBH VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=1.13999 scb=8.44443e-05 scc=9.17689e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=5.284 scb=0.00326881 scc=8.68818e-05
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@24 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=4.17894 scb=0.00212503
+ scc=8.30326e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=5.6e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@23 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=3.6279 scb=0.00186615
+ scc=8.2884e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@22 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.44e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@21 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.88e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@20 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@19 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@18 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@17 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@16 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@15 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@14 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@13 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@12 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@11 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@10 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@9 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@8 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@7 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@6 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M2 XI0/XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=3.125e-06 AD=2.1875e-13 AS=3.75e-13 PD=3.265e-06 PS=6.49e-06 M=1 sca=3.09215
+ scb=0.00283651 scc=0.000132595 lpccnr=2.85e-07 covpccnr=0 wrxcnr=2.8125e-06
+ sa=1.2e-07 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@5 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M2@8 XI0/XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=3.125e-06 AD=2.1875e-13 AS=2.1875e-13 PD=3.265e-06 PS=3.265e-06 M=1
+ sca=3.09215 scb=0.00283651 scc=0.000132595 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=2.8125e-06 sa=5.6e-07 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@4 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/XI0/M2@7 XI0/XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=3.125e-06 AD=2.1875e-13 AS=2.1875e-13 PD=3.265e-06 PS=3.265e-06 M=1
+ sca=3.09215 scb=0.00283651 scc=0.000132595 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=2.8125e-06 sa=1e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@3 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=2.534 scb=0.00179678
+ scc=8.28784e-05 lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06
+ sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M2@6 XI0/XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=3.125e-06 AD=2.1875e-13 AS=3.75e-13 PD=3.265e-06 PS=6.49e-06 M=1
+ sca=3.09215 scb=0.00283651 scc=0.000132595 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=2.8125e-06 sa=1.44e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1N@2 XI0/XI0/XI0/XI0/N2N XI0/XI0/XI0/XI0/N1N152
+ XI0/XI0/XI0/XI0/N1 XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13
+ AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06
+ PS=1.024e-05 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M2@5 XI0/XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=3.125e-06 AD=2.1875e-13 AS=3.75e-13 PD=3.265e-06 PS=6.49e-06 M=1
+ sca=3.09215 scb=0.00283651 scc=0.000132595 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=2.8125e-06 sa=1.2e-07 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@24 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=5.6e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M2@4 XI0/XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=3.125e-06 AD=2.1875e-13 AS=2.1875e-13 PD=3.265e-06 PS=3.265e-06 M=1
+ sca=3.09215 scb=0.00283651 scc=0.000132595 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=2.8125e-06 sa=5.6e-07 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@23 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=1e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M2@3 XI0/XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=3.125e-06 AD=2.1875e-13 AS=2.1875e-13 PD=3.265e-06 PS=3.265e-06 M=1
+ sca=3.09215 scb=0.00283651 scc=0.000132595 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=2.8125e-06 sa=1e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@22 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.44e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M2@2 XI0/XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet
+ L=3e-07 W=3.125e-06 AD=2.1875e-13 AS=3.75e-13 PD=3.265e-06 PS=6.49e-06 M=1
+ sca=3.09215 scb=0.00283651 scc=0.000132595 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=2.8125e-06 sa=1.44e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@21 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.88e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@20 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@19 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@18 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@17 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@16 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@15 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@14 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@13 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@12 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@11 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@10 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@9 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@8 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@7 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1
+ nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@6 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@5 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=2.534 scb=0.00179678 scc=8.28784e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@4 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=3.6279 scb=0.00186615 scc=8.2884e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@3 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=3.5e-13 PD=5.14e-06
+ PS=5.14e-06 M=1 sca=4.17894 scb=0.00212503 scc=8.30326e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XI0/M1P@2 XI0/XI0/XI0/VBN XI0/VCM XI0/XI0/XI0/XI0/N1
+ XI0/XI0/XI0/XI0/N1 egpfet L=3e-07 W=5e-06 AD=3.5e-13 AS=6e-13 PD=5.14e-06
+ PS=1.024e-05 M=1 sca=5.284 scb=0.00326881 scc=8.68818e-05 lpccnr=2.85e-07
+ covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XIRTN/RR1 TXP XI0/XI0/CM VDDHA_TX opppcres 188.174 M=1 w=5e-06
+ l=1.435e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI0/XI0/XIRTN/RR2 TXP XI0/XI0/CM VDDHA_TX opppcres 188.174 M=1 w=5e-06
+ l=1.435e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI0/XI0/XIRTN/RR3 TXP XI0/XI0/CM VDDHA_TX opppcres 188.174 M=1 w=5e-06
+ l=1.435e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI0/XI0/XIRTN/RR4 TXP XI0/XI0/CM VDDHA_TX opppcres 188.174 M=1 w=5e-06
+ l=1.435e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XX287/X24/X35/X126/X3/D0_noxref X287/X24/X35/X126/X3/noxref_2591 XI0/XI0/XI0/N1
+ diodenwx  AREA=1.52601e-09 perim=0.0001613 sizedup=0
XXI0/XI0/XI0/M3N TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=1.023e-11 PD=2.494e-05 PS=4.493e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=4.65e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M3N@22 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@21 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@20 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@19 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@18 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@17 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@16 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@15 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@14 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@13 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@12 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@11 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@10 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@9 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@8 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@7 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@6 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@5 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@4 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@3 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3N@2 TXP XI0/XI0/NN3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=1.023e-11 PD=2.494e-05 PS=4.493e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=4.65e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M4N TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=1.023e-11 PD=2.494e-05 PS=4.493e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=4.65e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@22 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@21 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@20 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@19 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@18 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@17 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@16 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@15 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@14 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@13 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@12 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@11 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@10 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@9 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@8 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@7 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@6 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@5 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@4 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@3 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4N@2 TXP XI0/XI0/NN3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=1.023e-11 PD=2.494e-05 PS=4.493e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=4.65e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX287/X24/X35/X126/X5/D0_noxref VSSA_TX VDDHA_TX diodenwx  AREA=1.60692e-11
+ perim=1.752e-05 sizedup=0
XXI0/XI0/XI0/RR2 TXP XI0/XI0/XI0/N1N798 VDDHA_TX opppcres 968.268 M=1 w=2e-06
+ l=3.08e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI0/XI0/MC2 VSSA_TX XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=5e-06 W=5e-06
+ AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=2.17174 scb=0.00193499
+ scc=0.000107095 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.3e-07
+ sb=1.3e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC2@8 VSSA_TX XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=5e-06
+ W=5e-06 AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=0.442158
+ scb=1.43115e-05 scc=2.13593e-09 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MPD2 XI0/XI0/XI0/N1N798 XI0/XI0/ENBH VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1 sca=8.2713
+ scb=0.00782352 scc=0.000835577 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.8e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MPD2@2 XI0/XI0/XI0/N1N798 XI0/XI0/ENBH VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1 sca=8.2713
+ scb=0.00782352 scc=0.000835577 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.8e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC2@7 VSSA_TX XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=5e-06
+ W=5e-06 AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC2@6 VSSA_TX XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=5e-06
+ W=5e-06 AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=0.442158
+ scb=1.43115e-05 scc=2.13593e-09 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@23 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=1.14755
+ scb=0.000590218 scc=6.64827e-06 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@24 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@25 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=1.14755
+ scb=0.000590218 scc=6.64827e-06 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@26 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=8.4e-13 AS=4.9e-13 PD=1.424e-05 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=5.6e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@2 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=1e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@3 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=1.44e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@4 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=1.88e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@5 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@6 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@7 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@8 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@9 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@10 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@11 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@12 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@13 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@14 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@15 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@16 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@17 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@18 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@19 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@20 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@21 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@22 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@23 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@24 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@25 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@26 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@27 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@28 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@29 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@30 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@31 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@32 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@33 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@34 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@35 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@36 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@37 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@38 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@39 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@40 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@41 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@42 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@43 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@44 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@45 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@46 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@47 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@48 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@49 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@50 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@51 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@52 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@53 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@54 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@55 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@56 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@57 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@58 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@59 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@60 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@61 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@62 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@63 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=8.4e-13 AS=4.9e-13 PD=1.424e-05 PS=7.14e-06 M=1
+ sca=0.274166 scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=1.5e-12 AS=8.75e-13 PD=2.524e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=5.6e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@2 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=1e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@3 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=1.44e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@4 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=1.88e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@5 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@6 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@7 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@8 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@9 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@10 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@11 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@12 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@13 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@14 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@15 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@16 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@17 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@18 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@19 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@20 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@21 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@22 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@23 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@24 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@25 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@26 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@27 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@28 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@29 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@30 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@31 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@32 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@33 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@34 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@35 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@36 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@37 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@38 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@39 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@40 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@41 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@42 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@43 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@44 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@45 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@46 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@47 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@48 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@49 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@50 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@51 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@52 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@53 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@54 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@55 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@56 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@57 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@58 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@59 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@60 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@61 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@62 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@63 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=1.5e-12 AS=8.75e-13 PD=2.524e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/XIRTP/RR1 TXN XI0/XI0/CM VDDHA_TX opppcres 188.174 M=1 w=5e-06
+ l=1.435e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI0/XI0/XIRTP/RR2 TXN XI0/XI0/CM VDDHA_TX opppcres 188.174 M=1 w=5e-06
+ l=1.435e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI0/XI0/XIRTP/RR3 TXN XI0/XI0/CM VDDHA_TX opppcres 188.174 M=1 w=5e-06
+ l=1.435e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI0/XI0/XIRTP/RR4 TXN XI0/XI0/CM VDDHA_TX opppcres 188.174 M=1 w=5e-06
+ l=1.435e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XX287/X24/X35/X127/X3/D0_noxref X287/X24/X35/X127/X3/noxref_2591 XI0/XI0/XI0/N1
+ diodenwx  AREA=1.52601e-09 perim=0.0001613 sizedup=0
XXI0/XI0/XI0/M3P TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=1.023e-11 PD=2.494e-05 PS=4.493e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=4.65e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M3P@22 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@21 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@20 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@19 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@18 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@17 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@16 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@15 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@14 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@13 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@12 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@11 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@10 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@9 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@8 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@7 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@6 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@5 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@4 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@3 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M3P@2 TXN XI0/XI0/NP3A XI0/XI0/XI0/N1 XI0/XI0/XI0/N1 egpfet
+ L=1.5e-07 W=2.2e-05 AD=3.234e-11 AS=1.023e-11 PD=2.494e-05 PS=4.493e-05 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06
+ sb=4.65e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M4P TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=1.023e-11 PD=2.494e-05 PS=4.493e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=4.65e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@22 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@21 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@20 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@19 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@18 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@17 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@16 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@15 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@14 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@13 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@12 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@11 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@10 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@9 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@8 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@7 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@6 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@5 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@4 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@3 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=9.24e-12 PD=2.494e-05 PS=2.284e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI0/M4P@2 TXN XI0/XI0/NP3B XI0/XI0/XI0/N2 VSSA_TX egnfet L=1.5e-07
+ W=2.2e-05 AD=3.234e-11 AS=1.023e-11 PD=2.494e-05 PS=4.493e-05 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.98e-05 sa=2.0083e-06 sb=4.65e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX287/X24/X35/X127/X5/D0_noxref VSSA_TX VDDHA_TX diodenwx  AREA=1.60692e-11
+ perim=1.752e-05 sizedup=0
XXI0/XI0/XI0/RR1 TXN XI0/XI0/XI0/N1N789 VDDHA_TX opppcres 968.268 M=1 w=2e-06
+ l=3.08e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI0/XI0/XI0/MC2@5 VSSA_TX XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=5e-06
+ W=5e-06 AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=2.17174
+ scb=0.00193499 scc=0.000107095 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC2@4 VSSA_TX XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=5e-06
+ W=5e-06 AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=0.442158
+ scb=1.43115e-05 scc=2.13593e-09 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MPD1 XI0/XI0/XI0/N1N789 XI0/XI0/ENBH VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1 sca=8.2713
+ scb=0.00782352 scc=0.000835577 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.8e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MPD1@2 XI0/XI0/XI0/N1N789 XI0/XI0/ENBH VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1 sca=8.2713
+ scb=0.00782352 scc=0.000835577 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.8e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC2@3 VSSA_TX XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=5e-06
+ W=5e-06 AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC2@2 VSSA_TX XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=5e-06
+ W=5e-06 AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=0.442158
+ scb=1.43115e-05 scc=2.13593e-09 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@27 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=1.14755
+ scb=0.000590218 scc=6.64827e-06 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@28 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@29 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=1.14755
+ scb=0.000590218 scc=6.64827e-06 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/MC1@30 VDDHA_TX XI0/VBP VDDHA_TX VDDHA_TX egpfet L=5e-06 W=5e-06
+ AD=6.5e-13 AS=6.5e-13 PD=1.026e-05 PS=1.026e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.3e-07 sb=1.3e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2P@64 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=8.4e-13 AS=4.9e-13 PD=1.424e-05 PS=7.14e-06 M=1
+ sca=0.274166 scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@2 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=5.6e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@3 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=1e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@4 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=1.44e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@5 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=1.88e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@6 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@7 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@8 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@9 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet L=3e-07
+ W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@10 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@11 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@12 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@13 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@14 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@15 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@16 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@17 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@18 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@19 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@20 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@21 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@22 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@23 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@24 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@25 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@26 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@27 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@28 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@29 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@30 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@31 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@32 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@33 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@34 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@35 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@36 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@37 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@38 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@39 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@40 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@41 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@42 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@43 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@44 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@45 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@46 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@47 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@48 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@49 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@50 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@51 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@52 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@53 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@54 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@55 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@56 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@57 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@58 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@59 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@60 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@61 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@62 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@63 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1 sca=0.274166
+ scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M2N@64 XI0/XI0/XI0/N2 XI0/XI0/XI0/VBN VSSA_TX VSSA_TX egnfet
+ L=3e-07 W=7e-06 AD=8.4e-13 AS=4.9e-13 PD=1.424e-05 PS=7.14e-06 M=1
+ sca=0.274166 scb=2.38475e-06 scc=7.10589e-11 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1P@64 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=1.5e-12 AS=8.75e-13 PD=2.524e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@2 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=5.6e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@3 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=1e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@4 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=1.44e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@5 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=1.88e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@6 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@7 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@8 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@9 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@10 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@11 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@12 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@13 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@14 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@15 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@16 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@17 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@18 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@19 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@20 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@21 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@22 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@23 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@24 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@25 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@26 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@27 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@28 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@29 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@30 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@31 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@32 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@33 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@34 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@35 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@36 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@37 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@38 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@39 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@40 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@41 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@42 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@43 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@44 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@45 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@46 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@47 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@48 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@49 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@50 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@51 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@52 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@53 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@54 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@55 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@56 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@57 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@58 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@59 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@60 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=1.88e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@61 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@62 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@63 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=8.75e-13 AS=8.75e-13 PD=1.264e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI0/M1N@64 XI0/XI0/XI0/N1 XI0/VBP VDDHA_TX VDDHA_TX egpfet L=3e-07
+ W=1.25e-05 AD=1.5e-12 AS=8.75e-13 PD=2.524e-05 PS=1.264e-05 M=1 sca=0.579718
+ scb=0.00033211 scc=5.73645e-06 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.125e-05
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XX287/X24/X36/D0_noxref VSS VDDHA_TX diodenwx  AREA=3.34642e-11 perim=2.386e-05
+ sizedup=0
XXI0/XI0/XI1/M9 XI0/XI0/NN3A XI0/XI0/XI1/S1 XI0/XI0/NN3B VSSA_TX egnfet
+ L=1.5e-07 W=2.5e-06 AD=3e-13 AS=1.75e-13 PD=5.24e-06 PS=2.64e-06 M=1
+ sca=0.640321 scb=2.00318e-05 scc=2.00916e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M9@4 XI0/XI0/NN3A XI0/XI0/XI1/S1 XI0/XI0/NN3B VSSA_TX egnfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1
+ sca=0.640321 scb=2.00318e-05 scc=2.00916e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M9@3 XI0/XI0/NN3A XI0/XI0/XI1/S1 XI0/XI0/NN3B VSSA_TX egnfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1
+ sca=0.640321 scb=2.00318e-05 scc=2.00916e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M9@2 XI0/XI0/NN3A XI0/XI0/XI1/S1 XI0/XI0/NN3B VSSA_TX egnfet
+ L=1.5e-07 W=2.5e-06 AD=3e-13 AS=1.75e-13 PD=5.24e-06 PS=2.64e-06 M=1
+ sca=0.640321 scb=2.00318e-05 scc=2.00916e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1 sca=1.1306
+ scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.8e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10@12 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10@12 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10@11 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10@11 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10@10 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=9.9e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10@10 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=9.9e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10@9 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.28e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10@9 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.28e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10@8 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.57e-06 sb=1.86e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10@8 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.57e-06 sb=1.86e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10@7 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.86e-06 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10@7 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.86e-06 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10@6 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10@6 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10@5 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10@5 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10@4 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10@4 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10@3 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10@3 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M10@2 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M10@2 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M8 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M8 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M8@6 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M8@6 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M8@5 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M8@5 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M8@4 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M8@4 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M8@3 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M8@3 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M8@2 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M8@2 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M6 XI0/XI0/XI1/XI0P/N1N28 XI0/XI0/XI1/XI0P/N1N29 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06
+ PS=3.24e-06 M=1 sca=1.31564 scb=0.000238286 scc=2.21595e-07 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.35e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M6 XI0/XI0/XI1/XI1P/N1N28 XI0/XI0/XI1/XI1P/N1N29 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06
+ PS=3.24e-06 M=1 sca=2.23358 scb=0.00029503 scc=2.31968e-07 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.35e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M6@2 XI0/XI0/XI1/XI0P/N1N28 XI0/XI0/XI1/XI0P/N1N29 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06
+ PS=3.24e-06 M=1 sca=1.31564 scb=0.000238286 scc=2.21595e-07 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.35e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M6@2 XI0/XI0/XI1/XI1P/N1N28 XI0/XI0/XI1/XI1P/N1N29 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06
+ PS=3.24e-06 M=1 sca=2.23358 scb=0.00029503 scc=2.31968e-07 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.35e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M4B XI0/XI0/XI1/XI0P/N1N50 VDDHA_TX VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1
+ sca=1.31564 scb=0.000238286 scc=2.21595e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.35e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M4B XI0/XI0/XI1/XI1P/N1N50 VSSA_TX VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1
+ sca=2.23358 scb=0.00029503 scc=2.31968e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.35e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M3B XI0/XI0/XI1/XI0P/N1N29 XI0/XI0/XI1/S1B
+ XI0/XI0/XI1/XI0P/N1N50 VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13
+ AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.31564 scb=0.000238286
+ scc=2.21595e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.35e-06 sa=4.1e-07 sb=7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI1P/M3B XI0/XI0/XI1/XI1P/N1N29 XI0/XI0/XI1/S1B
+ XI0/XI0/XI1/XI1P/N1N50 VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13
+ AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=2.23358 scb=0.00029503
+ scc=2.31968e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.35e-06 sa=4.1e-07 sb=7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI0P/M3A XI0/XI0/XI1/XI0P/N1N29 XI0/XI0/XI1/S1
+ XI0/XI0/XI1/XI0P/N1N42 VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13
+ AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.31564 scb=0.000238286
+ scc=2.21595e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.35e-06 sa=7e-07 sb=4.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI1P/M3A XI0/XI0/XI1/XI1P/N1N29 XI0/XI0/XI1/S1
+ XI0/XI0/XI1/XI1P/N1N42 VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13
+ AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=2.23358 scb=0.00029503
+ scc=2.31968e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.35e-06 sa=7e-07 sb=4.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI0P/M4A XI0/XI0/XI1/XI0P/N1N42 XI0/XI0/XI1/N1 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1
+ sca=1.31564 scb=0.000238286 scc=2.21595e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.35e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M4A XI0/XI0/XI1/XI1P/N1N42 XI0/XI0/XI1/N1 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1
+ sca=2.23358 scb=0.00029503 scc=2.31968e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.35e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M7 XI0/XI0/XI1/NN XI0/XI0/XI1/N1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=1.2e-13 PD=1.14e-06 PS=2.24e-06 M=1 sca=0.760516
+ scb=1.68732e-05 scc=5.36472e-10 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07
+ sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M7@6 XI0/XI0/XI1/NN XI0/XI0/XI1/N1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=7e-14 PD=1.14e-06 PS=1.14e-06 M=1 sca=0.760516
+ scb=1.68732e-05 scc=5.36472e-10 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07
+ sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M2 XI0/XI0/XI1/N1 XI0/XI0/NP2 XI0/XI0/XI1/NN VSSA_TX egnfet
+ L=1.5e-07 W=6e-07 AD=4.2e-14 AS=7.2e-14 PD=7.4e-07 PS=1.44e-06 M=1 sca=1.14059
+ scb=8.9985e-05 scc=1.25464e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.4e-07
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M7@5 XI0/XI0/XI1/NN XI0/XI0/XI1/N1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=7e-14 PD=1.14e-06 PS=1.14e-06 M=1 sca=0.760516
+ scb=1.68732e-05 scc=5.36472e-10 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07
+ sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M2@4 XI0/XI0/XI1/N1 XI0/XI0/NP2 XI0/XI0/XI1/NN VSSA_TX egnfet
+ L=1.5e-07 W=6e-07 AD=4.2e-14 AS=4.2e-14 PD=7.4e-07 PS=7.4e-07 M=1 sca=1.14059
+ scb=8.9985e-05 scc=1.25464e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.4e-07
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/X1I156/M2 XI0/XI0/XI1/N1N118 XI0/XI0/ENBH VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=1.14489 scb=8.59628e-05 scc=9.53026e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M7@4 XI0/XI0/XI1/NN XI0/XI0/XI1/N1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=7e-14 PD=1.14e-06 PS=1.14e-06 M=1 sca=0.760516
+ scb=1.68732e-05 scc=5.36472e-10 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07
+ sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M2@3 XI0/XI0/XI1/N1 XI0/XI0/NP2 XI0/XI0/XI1/NN VSSA_TX egnfet
+ L=1.5e-07 W=6e-07 AD=4.2e-14 AS=4.2e-14 PD=7.4e-07 PS=7.4e-07 M=1 sca=1.14059
+ scb=8.9985e-05 scc=1.25464e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.4e-07
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M7@3 XI0/XI0/XI1/NN XI0/XI0/XI1/N1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=7e-14 PD=1.14e-06 PS=1.14e-06 M=1 sca=0.760516
+ scb=1.68732e-05 scc=5.36472e-10 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07
+ sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M2@2 XI0/XI0/XI1/N1 XI0/XI0/NP2 XI0/XI0/XI1/NN VSSA_TX egnfet
+ L=1.5e-07 W=6e-07 AD=4.2e-14 AS=7.2e-14 PD=7.4e-07 PS=1.44e-06 M=1 sca=1.14059
+ scb=8.9985e-05 scc=1.25464e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.4e-07
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M7@2 XI0/XI0/XI1/NN XI0/XI0/XI1/N1 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=1.2e-13 PD=1.14e-06 PS=2.24e-06 M=1 sca=0.760516
+ scb=1.68732e-05 scc=5.36472e-10 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07
+ sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/X1I175/M2 XI0/XI0/XI1/S1B XI0/XI0/XI1/N1N118 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=1.14489
+ scb=8.59628e-05 scc=9.53026e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/X1I175/M2@2 XI0/XI0/XI1/S1B XI0/XI0/XI1/N1N118 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=4e-07 AD=2.8e-14 AS=2.8e-14 PD=5.4e-07 PS=5.4e-07 M=1
+ sca=1.14489 scb=8.59628e-05 scc=9.53026e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/X1I134/M2 XI0/XI0/XI1/S1 XI0/XI0/XI1/S1B VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=2.8e-14 PD=5.4e-07 PS=5.4e-07 M=1 sca=1.14489
+ scb=8.59628e-05 scc=9.53026e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/X1I134/M2@2 XI0/XI0/XI1/S1 XI0/XI0/XI1/S1B VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=1.14489
+ scb=8.59628e-05 scc=9.53026e-09 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M8 XI0/XI0/XI1/NN XI0/XI0/XI1/N2 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=1.2e-13 PD=1.14e-06 PS=2.24e-06 M=1 sca=0.760516
+ scb=1.68732e-05 scc=5.36472e-10 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07
+ sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M4 XI0/XI0/XI1/N2 XI0/XI0/NN2 XI0/XI0/XI1/NN VSSA_TX egnfet
+ L=1.5e-07 W=6e-07 AD=4.2e-14 AS=7.2e-14 PD=7.4e-07 PS=1.44e-06 M=1 sca=1.14059
+ scb=8.9985e-05 scc=1.25464e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.4e-07
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M8@6 XI0/XI0/XI1/NN XI0/XI0/XI1/N2 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=7e-14 PD=1.14e-06 PS=1.14e-06 M=1 sca=0.760516
+ scb=1.68732e-05 scc=5.36472e-10 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07
+ sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M4@4 XI0/XI0/XI1/N2 XI0/XI0/NN2 XI0/XI0/XI1/NN VSSA_TX egnfet
+ L=1.5e-07 W=6e-07 AD=4.2e-14 AS=4.2e-14 PD=7.4e-07 PS=7.4e-07 M=1 sca=1.14059
+ scb=8.9985e-05 scc=1.25464e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.4e-07
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M8@5 XI0/XI0/XI1/NN XI0/XI0/XI1/N2 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=7e-14 PD=1.14e-06 PS=1.14e-06 M=1 sca=0.760516
+ scb=1.68732e-05 scc=5.36472e-10 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07
+ sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M4@3 XI0/XI0/XI1/N2 XI0/XI0/NN2 XI0/XI0/XI1/NN VSSA_TX egnfet
+ L=1.5e-07 W=6e-07 AD=4.2e-14 AS=4.2e-14 PD=7.4e-07 PS=7.4e-07 M=1 sca=1.14059
+ scb=8.9985e-05 scc=1.25464e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.4e-07
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M8@4 XI0/XI0/XI1/NN XI0/XI0/XI1/N2 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=7e-14 PD=1.14e-06 PS=1.14e-06 M=1 sca=0.228155
+ scb=5.06196e-06 scc=1.60942e-10 lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07
+ sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M4@2 XI0/XI0/XI1/N2 XI0/XI0/NN2 XI0/XI0/XI1/NN VSSA_TX egnfet
+ L=1.5e-07 W=6e-07 AD=4.2e-14 AS=7.2e-14 PD=7.4e-07 PS=1.44e-06 M=1 sca=1.14059
+ scb=8.9985e-05 scc=1.25464e-08 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.4e-07
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M8@3 XI0/XI0/XI1/NN XI0/XI0/XI1/N2 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=7e-14 PD=1.14e-06 PS=1.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07 sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M8@2 XI0/XI0/XI1/NN XI0/XI0/XI1/N2 VSSA_TX VSSA_TX egnfet L=1.5e-07
+ W=1e-06 AD=7e-14 AS=1.2e-13 PD=1.14e-06 PS=2.24e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=9e-07 sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M4A XI0/XI0/XI1/XI1N/N1N42 XI0/XI0/XI1/N2 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1
+ sca=2.23358 scb=0.00029503 scc=2.31968e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.35e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M4A XI0/XI0/XI1/XI0N/N1N42 XI0/XI0/XI1/N2 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1
+ sca=1.31564 scb=0.000238286 scc=2.21595e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.35e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M3A XI0/XI0/XI1/XI1N/N1N29 XI0/XI0/XI1/S1
+ XI0/XI0/XI1/XI1N/N1N42 VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13
+ AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=2.23358 scb=0.00029503
+ scc=2.31968e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.35e-06 sa=4.1e-07 sb=7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI0N/M3A XI0/XI0/XI1/XI0N/N1N29 XI0/XI0/XI1/S1
+ XI0/XI0/XI1/XI0N/N1N42 VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13
+ AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.31564 scb=0.000238286
+ scc=2.21595e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.35e-06 sa=4.1e-07 sb=7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI1N/M3B XI0/XI0/XI1/XI1N/N1N29 XI0/XI0/XI1/S1B
+ XI0/XI0/XI1/XI1N/N1N50 VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13
+ AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=2.23358 scb=0.00029503
+ scc=2.31968e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.35e-06 sa=7e-07 sb=4.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI0N/M3B XI0/XI0/XI1/XI0N/N1N29 XI0/XI0/XI1/S1B
+ XI0/XI0/XI1/XI0N/N1N50 VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13
+ AS=1.05e-13 PD=1.64e-06 PS=1.64e-06 M=1 sca=1.31564 scb=0.000238286
+ scc=2.21595e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.35e-06 sa=7e-07 sb=4.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI1N/M4B XI0/XI0/XI1/XI1N/N1N50 VSSA_TX VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1
+ sca=2.23358 scb=0.00029503 scc=2.31968e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.35e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M4B XI0/XI0/XI1/XI0N/N1N50 VDDHA_TX VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06 PS=3.24e-06 M=1
+ sca=1.31564 scb=0.000238286 scc=2.21595e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.35e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M6 XI0/XI0/XI1/XI1N/N1N28 XI0/XI0/XI1/XI1N/N1N29 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06
+ PS=3.24e-06 M=1 sca=2.23358 scb=0.00029503 scc=2.31968e-07 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.35e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M6 XI0/XI0/XI1/XI0N/N1N28 XI0/XI0/XI1/XI0N/N1N29 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06
+ PS=3.24e-06 M=1 sca=1.31564 scb=0.000238286 scc=2.21595e-07 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.35e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M6@2 XI0/XI0/XI1/XI1N/N1N28 XI0/XI0/XI1/XI1N/N1N29 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06
+ PS=3.24e-06 M=1 sca=2.23358 scb=0.00029503 scc=2.31968e-07 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.35e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M6@2 XI0/XI0/XI1/XI0N/N1N28 XI0/XI0/XI1/XI0N/N1N29 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=1.5e-06 AD=1.05e-13 AS=1.8e-13 PD=1.64e-06
+ PS=3.24e-06 M=1 sca=1.31564 scb=0.000238286 scc=2.21595e-07 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=1.35e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M8 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M8 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M8@6 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M8@6 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M8@5 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M8@5 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M8@4 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M8@4 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M8@3 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M8@3 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M8@2 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06
+ M=1 sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M8@2 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VSSA_TX
+ VSSA_TX egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06
+ M=1 sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX egnfet
+ L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1 sca=1.1306
+ scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.8e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10@12 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10@12 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=4.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10@11 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10@11 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10@10 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=9.9e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10@10 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=9.9e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10@9 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.28e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10@9 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.28e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10@8 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.57e-06 sb=1.86e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10@8 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.57e-06 sb=1.86e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10@7 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.86e-06 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10@7 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=1.86e-06 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10@6 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10@6 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10@5 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10@5 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10@4 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10@4 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10@3 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10@3 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=1.4e-13 PD=2.14e-06 PS=2.14e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M10@2 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1
+ sca=2.36183 scb=0.000423719 scc=4.89349e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M10@2 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VSSA_TX VSSA_TX
+ egnfet L=1.5e-07 W=2e-06 AD=1.4e-13 AS=2.4e-13 PD=2.14e-06 PS=4.24e-06 M=1
+ sca=1.1306 scb=0.000179402 scc=1.66198e-07 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.8e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M11 XI0/XI0/NP3A XI0/XI0/XI1/S1 XI0/XI0/NP3B VSSA_TX egnfet
+ L=1.5e-07 W=2.5e-06 AD=3e-13 AS=1.75e-13 PD=5.24e-06 PS=2.64e-06 M=1
+ sca=0.640321 scb=2.00318e-05 scc=2.00916e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M11@4 XI0/XI0/NP3A XI0/XI0/XI1/S1 XI0/XI0/NP3B VSSA_TX egnfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1
+ sca=0.640321 scb=2.00318e-05 scc=2.00916e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M11@3 XI0/XI0/NP3A XI0/XI0/XI1/S1 XI0/XI0/NP3B VSSA_TX egnfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1
+ sca=0.640321 scb=2.00318e-05 scc=2.00916e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M11@2 XI0/XI0/NP3A XI0/XI0/XI1/S1 XI0/XI0/NP3B VSSA_TX egnfet
+ L=1.5e-07 W=2.5e-06 AD=3e-13 AS=1.75e-13 PD=5.24e-06 PS=2.64e-06 M=1
+ sca=0.640321 scb=2.00318e-05 scc=2.00916e-09 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M10 XI0/XI0/NN3B XI0/XI0/XI1/S1B XI0/XI0/NN3A VDDHA_TX egpfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1
+ sca=5.2516 scb=0.00349131 scc=9.22571e-05 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M10@4 XI0/XI0/NN3B XI0/XI0/XI1/S1B XI0/XI0/NN3A VDDHA_TX egpfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1
+ sca=4.67477 scb=0.00302297 scc=9.1528e-05 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M10@3 XI0/XI0/NN3B XI0/XI0/XI1/S1B XI0/XI0/NN3A VDDHA_TX egpfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1
+ sca=4.30317 scb=0.00284904 scc=9.14438e-05 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M10@2 XI0/XI0/NN3B XI0/XI0/XI1/S1B XI0/XI0/NN3A VDDHA_TX egpfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1
+ sca=3.11007 scb=0.00275157 scc=9.14331e-05 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06 PS=1.424e-05 M=1
+ sca=3.13 scb=0.002644 scc=0.000131154 lpccnr=1.5e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06 PS=1.424e-05 M=1
+ sca=5.62279 scb=0.00379772 scc=0.000133358 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9@12 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.12068 scb=0.00263455 scc=0.000131129 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=4.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9@12 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=4.89734 scb=0.00306314 scc=0.000131386 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=4.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9@11 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.11486 scb=0.00263099 scc=0.000131126 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9@11 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=4.44498 scb=0.00278632 scc=0.000131155 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9@10 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.11099 scb=0.00262969 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=9.9e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9@10 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=4.14402 scb=0.00268496 scc=0.000131129 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=9.9e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9@9 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.28e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9@9 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.28e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9@8 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.57e-06 sb=1.86e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9@8 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.57e-06 sb=1.86e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M1B XI0/XI0/XI1/XI0P/N1N52 VDDHA_TX VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06 PS=1.074e-05 M=1
+ sca=2.57335 scb=0.0019486 scc=0.000109028 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=4.725e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M1B XI0/XI0/XI1/XI1P/N1N52 VSSA_TX VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06 PS=1.074e-05 M=1
+ sca=4.32859 scb=0.00237201 scc=0.000109282 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=4.725e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M2B XI0/XI0/XI1/XI0P/N1N29 XI0/XI0/XI1/S1
+ XI0/XI0/XI1/XI0P/N1N52 VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13
+ AS=3.675e-13 PD=5.39e-06 PS=5.39e-06 M=1 sca=2.59132 scb=0.00196679
+ scc=0.000109077 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.725e-06 sa=4.1e-07 sb=7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI1P/M2B XI0/XI0/XI1/XI1P/N1N29 XI0/XI0/XI1/S1
+ XI0/XI0/XI1/XI1P/N1N52 VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13
+ AS=3.675e-13 PD=5.39e-06 PS=5.39e-06 M=1 sca=5.05404 scb=0.00310659
+ scc=0.000111255 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.725e-06 sa=4.1e-07 sb=7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI0P/M2A XI0/XI0/XI1/XI0P/N1N29 XI0/XI0/XI1/S1B
+ XI0/XI0/XI1/XI0P/N1N38 VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13
+ AS=3.675e-13 PD=5.39e-06 PS=5.39e-06 M=1 sca=2.62283 scb=0.00201308
+ scc=0.00010948 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.725e-06 sa=7e-07 sb=4.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI1P/M2A XI0/XI0/XI1/XI1P/N1N29 XI0/XI0/XI1/S1B
+ XI0/XI0/XI1/XI1P/N1N38 VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13
+ AS=3.675e-13 PD=5.39e-06 PS=5.39e-06 M=1 sca=6.32679 scb=0.00497633
+ scc=0.000127523 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.725e-06 sa=7e-07 sb=4.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI0P/M1A XI0/XI0/XI1/XI0P/N1N38 XI0/XI0/XI1/N1 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06 PS=1.074e-05
+ M=1 sca=2.686 scb=0.00212337 scc=0.000112619 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=4.725e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M1A XI0/XI0/XI1/XI1P/N1N38 XI0/XI0/XI1/N1 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06 PS=1.074e-05
+ M=1 sca=8.87783 scb=0.00943022 scc=0.000254303 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=4.725e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M5 XI0/XI0/XI1/NP XI0/XI0/XI1/N1 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=3e-06 AD=2.1e-13 AS=3.6e-13 PD=3.14e-06 PS=6.24e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M5@6 XI0/XI0/XI1/NP XI0/XI0/XI1/N1 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=3e-06 AD=2.1e-13 AS=2.1e-13 PD=3.14e-06 PS=3.14e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M5@5 XI0/XI0/XI1/NP XI0/XI0/XI1/N1 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=3e-06 AD=2.1e-13 AS=2.1e-13 PD=3.14e-06 PS=3.14e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M5@4 XI0/XI0/XI1/NP XI0/XI0/XI1/N1 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=3e-06 AD=2.1e-13 AS=2.1e-13 PD=3.14e-06 PS=3.14e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M5@3 XI0/XI0/XI1/NP XI0/XI0/XI1/N1 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=3e-06 AD=2.1e-13 AS=2.1e-13 PD=3.14e-06 PS=3.14e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M1 XI0/XI0/XI1/N1 XI0/XI0/NP2 XI0/XI0/XI1/NP VDDHA_TX egpfet
+ L=1.5e-07 W=2.1e-06 AD=1.47e-13 AS=2.52e-13 PD=2.24e-06 PS=4.44e-06 M=1
+ sca=3.5641 scb=0.00327377 scc=0.000108849 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.89e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M5@2 XI0/XI0/XI1/NP XI0/XI0/XI1/N1 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=3e-06 AD=2.1e-13 AS=3.6e-13 PD=3.14e-06 PS=6.24e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M1@4 XI0/XI0/XI1/N1 XI0/XI0/NP2 XI0/XI0/XI1/NP VDDHA_TX egpfet
+ L=1.5e-07 W=2.1e-06 AD=1.47e-13 AS=1.47e-13 PD=2.24e-06 PS=2.24e-06 M=1
+ sca=3.5641 scb=0.00327377 scc=0.000108849 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.89e-06 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/X1I156/M1 XI0/XI0/XI1/N1N118 XI0/XI0/ENBH VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1
+ sca=12.3736 scb=0.0141021 scc=0.000457256 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.26e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M1@3 XI0/XI0/XI1/N1 XI0/XI0/NP2 XI0/XI0/XI1/NP VDDHA_TX egpfet
+ L=1.5e-07 W=2.1e-06 AD=1.47e-13 AS=1.47e-13 PD=2.24e-06 PS=2.24e-06 M=1
+ sca=3.5641 scb=0.00327377 scc=0.000108849 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.89e-06 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M1@2 XI0/XI0/XI1/N1 XI0/XI0/NP2 XI0/XI0/XI1/NP VDDHA_TX egpfet
+ L=1.5e-07 W=2.1e-06 AD=1.47e-13 AS=2.52e-13 PD=2.24e-06 PS=4.44e-06 M=1
+ sca=3.5641 scb=0.00327377 scc=0.000108849 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.89e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/X1I175/M1 XI0/XI0/XI1/S1B XI0/XI0/XI1/N1N118 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06 PS=3.04e-06 M=1
+ sca=8.31129 scb=0.00650978 scc=0.000296 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.26e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/X1I175/M1@2 XI0/XI0/XI1/S1B XI0/XI0/XI1/N1N118 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=9.8e-14 PD=1.54e-06 PS=1.54e-06 M=1
+ sca=8.32841 scb=0.00652637 scc=0.000296011 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.26e-06 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/X1I134/M1 XI0/XI0/XI1/S1 XI0/XI0/XI1/S1B VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=9.8e-14 PD=1.54e-06 PS=1.54e-06 M=1
+ sca=7.75987 scb=0.0068106 scc=0.000296382 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.26e-06 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/X1I134/M1@2 XI0/XI0/XI1/S1 XI0/XI0/XI1/S1B VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06 PS=3.04e-06 M=1
+ sca=8.57539 scb=0.00772015 scc=0.000299559 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.26e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M3 XI0/XI0/XI1/N2 XI0/XI0/NN2 XI0/XI0/XI1/NP VDDHA_TX egpfet
+ L=1.5e-07 W=2.1e-06 AD=1.47e-13 AS=2.52e-13 PD=2.24e-06 PS=4.44e-06 M=1
+ sca=3.5641 scb=0.00327377 scc=0.000108849 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.89e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M3@4 XI0/XI0/XI1/N2 XI0/XI0/NN2 XI0/XI0/XI1/NP VDDHA_TX egpfet
+ L=1.5e-07 W=2.1e-06 AD=1.47e-13 AS=1.47e-13 PD=2.24e-06 PS=2.24e-06 M=1
+ sca=3.5641 scb=0.00327377 scc=0.000108849 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.89e-06 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M3@3 XI0/XI0/XI1/N2 XI0/XI0/NN2 XI0/XI0/XI1/NP VDDHA_TX egpfet
+ L=1.5e-07 W=2.1e-06 AD=1.47e-13 AS=1.47e-13 PD=2.24e-06 PS=2.24e-06 M=1
+ sca=3.5641 scb=0.00327377 scc=0.000108849 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.89e-06 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M6 XI0/XI0/XI1/NP XI0/XI0/XI1/N2 VDDHA_TX VDDHA_TX egpfet L=1.5e-07
+ W=3e-06 AD=2.1e-13 AS=3.6e-13 PD=3.14e-06 PS=6.24e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M3@2 XI0/XI0/XI1/N2 XI0/XI0/NN2 XI0/XI0/XI1/NP VDDHA_TX egpfet
+ L=1.5e-07 W=2.1e-06 AD=1.47e-13 AS=2.52e-13 PD=2.24e-06 PS=4.44e-06 M=1
+ sca=3.5641 scb=0.00327377 scc=0.000108849 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=1.89e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M6@6 XI0/XI0/XI1/NP XI0/XI0/XI1/N2 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=3e-06 AD=2.1e-13 AS=2.1e-13 PD=3.14e-06 PS=3.14e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M6@5 XI0/XI0/XI1/NP XI0/XI0/XI1/N2 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=3e-06 AD=2.1e-13 AS=2.1e-13 PD=3.14e-06 PS=3.14e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M6@4 XI0/XI0/XI1/NP XI0/XI0/XI1/N2 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=3e-06 AD=2.1e-13 AS=2.1e-13 PD=3.14e-06 PS=3.14e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M6@3 XI0/XI0/XI1/NP XI0/XI0/XI1/N2 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=3e-06 AD=2.1e-13 AS=2.1e-13 PD=3.14e-06 PS=3.14e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M6@2 XI0/XI0/XI1/NP XI0/XI0/XI1/N2 VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=3e-06 AD=2.1e-13 AS=3.6e-13 PD=3.14e-06 PS=6.24e-06 M=1 sca=1.5625
+ scb=0.000763136 scc=6.28992e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.7e-06
+ sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M1A XI0/XI0/XI1/XI1N/N1N38 XI0/XI0/XI1/N2 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06 PS=1.074e-05
+ M=1 sca=8.87783 scb=0.00943022 scc=0.000254303 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=4.725e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M1A XI0/XI0/XI1/XI0N/N1N38 XI0/XI0/XI1/N2 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06 PS=1.074e-05
+ M=1 sca=2.686 scb=0.00212337 scc=0.000112619 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=4.725e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M2A XI0/XI0/XI1/XI1N/N1N29 XI0/XI0/XI1/S1B
+ XI0/XI0/XI1/XI1N/N1N38 VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13
+ AS=3.675e-13 PD=5.39e-06 PS=5.39e-06 M=1 sca=6.32679 scb=0.00497633
+ scc=0.000127523 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.725e-06 sa=4.1e-07 sb=7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI0N/M2A XI0/XI0/XI1/XI0N/N1N29 XI0/XI0/XI1/S1B
+ XI0/XI0/XI1/XI0N/N1N38 VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13
+ AS=3.675e-13 PD=5.39e-06 PS=5.39e-06 M=1 sca=2.62283 scb=0.00201308
+ scc=0.00010948 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.725e-06 sa=4.1e-07 sb=7e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI1N/M2B XI0/XI0/XI1/XI1N/N1N29 XI0/XI0/XI1/S1
+ XI0/XI0/XI1/XI1N/N1N52 VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13
+ AS=3.675e-13 PD=5.39e-06 PS=5.39e-06 M=1 sca=5.05404 scb=0.00310659
+ scc=0.000111255 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.725e-06 sa=7e-07 sb=4.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI0N/M2B XI0/XI0/XI1/XI0N/N1N29 XI0/XI0/XI1/S1
+ XI0/XI0/XI1/XI0N/N1N52 VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13
+ AS=3.675e-13 PD=5.39e-06 PS=5.39e-06 M=1 sca=2.59132 scb=0.00196679
+ scc=0.000109077 lpccnr=1.5e-07 covpccnr=0 wrxcnr=4.725e-06 sa=7e-07 sb=4.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI0/XI0/XI1/XI1N/M1B XI0/XI0/XI1/XI1N/N1N52 VSSA_TX VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06 PS=1.074e-05 M=1
+ sca=4.32859 scb=0.00237201 scc=0.000109282 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=4.725e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M1B XI0/XI0/XI1/XI0N/N1N52 VDDHA_TX VDDHA_TX VDDHA_TX egpfet
+ L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06 PS=1.074e-05 M=1
+ sca=2.57335 scb=0.0019486 scc=0.000109028 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=4.725e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.86e-06 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.86e-06 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9@12 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=2.0083e-06 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9@12 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=2.0083e-06 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9@11 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=4.14402 scb=0.00268496 scc=0.000131129 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=2.0083e-06 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9@11 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.11099 scb=0.00262969 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=2.0083e-06 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9@10 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=4.44498 scb=0.00278632 scc=0.000131155 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=2.0083e-06 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9@10 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.11486 scb=0.00263099 scc=0.000131126 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=2.0083e-06 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9@9 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=4.89734 scb=0.00306314 scc=0.000131386 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=2.0083e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9@9 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.12068 scb=0.00263455 scc=0.000131129 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=2.0083e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9@8 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06 PS=1.424e-05 M=1
+ sca=5.62279 scb=0.00379772 scc=0.000133358 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9@8 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06 PS=1.424e-05 M=1
+ sca=3.13 scb=0.002644 scc=0.000131154 lpccnr=1.5e-07 covpccnr=0 wrxcnr=6.3e-06
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M12 XI0/XI0/NP3B XI0/XI0/XI1/S1B XI0/XI0/NP3A VDDHA_TX egpfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1
+ sca=3.11007 scb=0.00275157 scc=9.14331e-05 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M12@4 XI0/XI0/NP3B XI0/XI0/XI1/S1B XI0/XI0/NP3A VDDHA_TX egpfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1
+ sca=4.30317 scb=0.00284904 scc=9.14438e-05 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M12@3 XI0/XI0/NP3B XI0/XI0/XI1/S1B XI0/XI0/NP3A VDDHA_TX egpfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=1.75e-13 PD=2.64e-06 PS=2.64e-06 M=1
+ sca=4.67477 scb=0.00302297 scc=9.1528e-05 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/M12@2 XI0/XI0/NP3B XI0/XI0/XI1/S1B XI0/XI0/NP3A VDDHA_TX egpfet
+ L=1.5e-07 W=2.5e-06 AD=1.75e-13 AS=3e-13 PD=2.64e-06 PS=5.24e-06 M=1
+ sca=5.2516 scb=0.00349131 scc=9.22571e-05 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.25e-06 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XX287/X24/X36/X209/D0_noxref VSS VDDHA_TX diodenwx  AREA=1.08528e-10
+ perim=4.303e-05 sizedup=0
XXI0/XI0/XI1/XI1P/M5 XI0/XI0/XI1/XI1P/N1N28 XI0/XI0/XI1/XI1P/N1N29 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06
+ PS=1.074e-05 M=1 sca=2.52879 scb=0.00193785 scc=0.000109022 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=4.725e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M5@2 XI0/XI0/XI1/XI1P/N1N28 XI0/XI0/XI1/XI1P/N1N29 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06
+ PS=1.074e-05 M=1 sca=2.52879 scb=0.00193785 scc=0.000109022 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=4.725e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M7 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06
+ PS=1.424e-05 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M7@6 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M7@5 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M7@4 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M7@3 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M7@2 XI0/XI0/XI1/XI1P/N1N25 XI0/XI0/XI1/XI1P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06
+ PS=1.424e-05 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9@7 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06 PS=1.424e-05 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9@6 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=4.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9@5 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9@4 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=9.9e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9@3 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.28e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1P/M9@2 XI0/XI0/NN3B XI0/XI0/XI1/XI1P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.57e-06 sb=1.86e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M5 XI0/XI0/XI1/XI0P/N1N28 XI0/XI0/XI1/XI0P/N1N29 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06
+ PS=1.074e-05 M=1 sca=2.52879 scb=0.00193785 scc=0.000109022 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=4.725e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M5@2 XI0/XI0/XI1/XI0P/N1N28 XI0/XI0/XI1/XI0P/N1N29 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06
+ PS=1.074e-05 M=1 sca=2.52879 scb=0.00193785 scc=0.000109022 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=4.725e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M7 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06
+ PS=1.424e-05 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M7@6 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M7@5 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M7@4 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M7@3 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M7@2 XI0/XI0/XI1/XI0P/N1N25 XI0/XI0/XI1/XI0P/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06
+ PS=1.424e-05 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9@7 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06 PS=1.424e-05 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9@6 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=4.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9@5 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9@4 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=9.9e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9@3 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.28e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0P/M9@2 XI0/XI0/NN3A XI0/XI0/XI1/XI0P/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.57e-06 sb=1.86e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XX287/X24/X36/X210/D0_noxref VSS VDDHA_TX diodenwx  AREA=1.08528e-10
+ perim=4.303e-05 sizedup=0
XXI0/XI0/XI1/XI1N/M5 XI0/XI0/XI1/XI1N/N1N28 XI0/XI0/XI1/XI1N/N1N29 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06
+ PS=1.074e-05 M=1 sca=2.52879 scb=0.00193785 scc=0.000109022 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=4.725e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M5@2 XI0/XI0/XI1/XI1N/N1N28 XI0/XI0/XI1/XI1N/N1N29 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06
+ PS=1.074e-05 M=1 sca=2.52879 scb=0.00193785 scc=0.000109022 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=4.725e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M7 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06
+ PS=1.424e-05 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M7@6 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M7@5 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M7@4 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M7@3 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M7@2 XI0/XI0/XI1/XI1N/N1N25 XI0/XI0/XI1/XI1N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06
+ PS=1.424e-05 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9@7 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06 PS=1.424e-05 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9@6 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=4.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9@5 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9@4 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=9.9e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9@3 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.28e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI1N/M9@2 XI0/XI0/NP3B XI0/XI0/XI1/XI1N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.57e-06 sb=1.86e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M5 XI0/XI0/XI1/XI0N/N1N28 XI0/XI0/XI1/XI0N/N1N29 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06
+ PS=1.074e-05 M=1 sca=2.52879 scb=0.00193785 scc=0.000109022 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=4.725e-06 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M5@2 XI0/XI0/XI1/XI0N/N1N28 XI0/XI0/XI1/XI0N/N1N29 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=5.25e-06 AD=3.675e-13 AS=6.3e-13 PD=5.39e-06
+ PS=1.074e-05 M=1 sca=2.52879 scb=0.00193785 scc=0.000109022 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=4.725e-06 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M7 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06
+ PS=1.424e-05 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.2e-07 sb=1.57e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M7@6 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=4.1e-07 sb=1.28e-06 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M7@5 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=7e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M7@4 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=9.9e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M7@3 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06
+ PS=7.14e-06 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.28e-06 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M7@2 XI0/XI0/XI1/XI0N/N1N25 XI0/XI0/XI1/XI0N/N1N28 VDDHA_TX
+ VDDHA_TX egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06
+ PS=1.424e-05 M=1 sca=3.10159 scb=0.00263164 scc=0.000132025 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=6.3e-06 sa=1.57e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9@7 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=8.4e-13 PD=7.14e-06 PS=1.424e-05 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9@6 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=4.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9@5 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=7e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9@4 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=9.9e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9@3 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.28e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI0/XI0/XI1/XI0N/M9@2 XI0/XI0/NP3A XI0/XI0/XI1/XI0N/N1N25 VDDHA_TX VDDHA_TX
+ egpfet L=1.5e-07 W=7e-06 AD=4.9e-13 AS=4.9e-13 PD=7.14e-06 PS=7.14e-06 M=1
+ sca=3.09753 scb=0.00262897 scc=0.000131125 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=6.3e-06 sa=1.57e-06 sb=1.86e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@512 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@511 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@510 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@509 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@508 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@507 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@506 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@505 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@504 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=5.25548 scb=0.0046872
+ scc=0.000346407 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@503 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@502 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@501 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@500 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@499 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@498 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@497 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@496 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@495 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@494 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@493 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@492 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@491 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@490 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@489 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@488 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@487 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@486 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@485 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@484 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@483 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@482 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@481 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@480 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@479 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@478 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@477 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@476 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@475 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@474 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@473 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@472 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@471 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@470 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@469 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@468 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@467 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@466 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@465 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@464 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@463 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@462 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@461 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@460 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@459 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@458 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=5.3309 scb=0.00475363
+ scc=0.000349818 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@457 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@456 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@455 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@454 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@453 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@452 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@451 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@450 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@449 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@448 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@447 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@446 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@445 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@444 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@443 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@442 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@441 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@440 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@439 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@438 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@437 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@436 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@435 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@434 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@433 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@432 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@431 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@430 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@429 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@428 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@427 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@426 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@425 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@424 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@423 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@422 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@421 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@420 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@419 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@418 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@417 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@416 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@415 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@414 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@413 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@412 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@411 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@410 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@409 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@408 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@407 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@406 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@405 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@404 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@403 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@402 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@401 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@400 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@399 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@398 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@397 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@396 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@395 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@394 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@393 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@392 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@391 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@390 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@389 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@388 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@387 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@386 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@385 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@384 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@383 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@382 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@381 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@380 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@379 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@378 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@377 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@376 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@375 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@374 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@373 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@372 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@371 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@370 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@369 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@368 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@367 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@366 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@365 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@364 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@363 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@362 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@361 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@360 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@359 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@358 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@357 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@356 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@355 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@354 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@353 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@352 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@351 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@350 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@349 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@348 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@347 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@346 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@345 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@344 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@343 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@342 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@341 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@340 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@339 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@338 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@337 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@336 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@335 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@334 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@333 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@332 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@331 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@330 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@329 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@328 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@327 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@326 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@325 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@324 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@323 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@322 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@321 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@320 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@319 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@318 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@317 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@316 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@315 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@314 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@313 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@312 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@311 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@310 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@309 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@308 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@307 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@306 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@305 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@304 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@303 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@302 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@301 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@300 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@299 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@298 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@297 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@296 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@295 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@294 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@293 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@292 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@291 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@290 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@289 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@288 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@287 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@286 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@285 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@284 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@283 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@282 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@281 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@280 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@279 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@278 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@277 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@276 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@275 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@274 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@273 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@272 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@271 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@270 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@269 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@268 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@267 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@266 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@265 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@264 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@263 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@262 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@261 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@260 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@259 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@258 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@257 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@256 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@255 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@254 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@253 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@252 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@251 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@250 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@249 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@248 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@247 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@246 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@245 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@244 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@243 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@242 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@241 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@240 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@239 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@238 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@237 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@236 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@235 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@234 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@233 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@232 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@231 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@230 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@229 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@228 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@227 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@226 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@225 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@224 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@223 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@222 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@221 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@220 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@219 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@218 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@217 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@216 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@215 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@214 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@213 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@212 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@211 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@210 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@209 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@208 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@207 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@206 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@205 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@204 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@203 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@202 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@201 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@200 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@199 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@198 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@197 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@196 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@195 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@194 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@193 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@192 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@191 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@190 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@189 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@188 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@187 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@186 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@185 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@184 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@183 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@182 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@181 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@180 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@179 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@178 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@177 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@176 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@175 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@174 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@173 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@172 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@171 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@170 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@169 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@168 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@167 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@166 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@165 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@164 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@163 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@162 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@161 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@160 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@159 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@158 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@157 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@156 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@155 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@154 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@153 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@152 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@151 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@150 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@149 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15255 scb=0.00189618
+ scc=9.73738e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@148 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@147 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@146 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@145 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=5.25548 scb=0.0046872
+ scc=0.000346407 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@144 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@143 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@142 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@141 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@140 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@139 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@138 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@137 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@136 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@135 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@134 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@133 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@132 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@131 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@130 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@129 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@128 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@127 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@126 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@125 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@124 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@123 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@122 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@121 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@120 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@119 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@118 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@117 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@116 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@115 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@114 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@113 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@112 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@111 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@110 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@109 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@108 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@107 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@106 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@105 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@104 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@103 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@102 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@101 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@100 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@99 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@98 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@97 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@96 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@95 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@94 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@93 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0.417892 scb=1.03815e-05
+ scc=1.08339e-09 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@92 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@91 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@90 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@89 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@88 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@87 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@86 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@85 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@84 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@83 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@82 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@81 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@80 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@79 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@78 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@77 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@76 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@75 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@74 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@73 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@72 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@71 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@70 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0.417892 scb=1.03815e-05
+ scc=1.08339e-09 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@69 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0.417892 scb=1.03815e-05
+ scc=1.08339e-09 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@68 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@67 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@66 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@65 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@64 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@63 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@62 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@61 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@60 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@59 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@58 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@57 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@56 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@55 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@54 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@53 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@52 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@51 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@50 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@49 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@48 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@47 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@46 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@45 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@44 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@43 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@42 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@41 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@40 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@39 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@38 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@37 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@36 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@35 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@34 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@33 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@32 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@31 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@30 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@29 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@28 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@27 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.504e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC1@26 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@25 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=3.2516 scb=0.00292199
+ scc=0.000255758 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@24 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.5726 scb=0.00190846
+ scc=9.74723e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@23 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@22 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@21 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@20 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@19 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@18 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@17 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@16 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@15 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@14 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@13 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@12 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@11 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@10 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@9 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@8 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@7 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@6 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@5 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@4 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@3 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC1@2 VDDHA_TX VSSA_TX VDDHA_TX VDDHA_TX pfet L=5e-06 W=5e-06 AD=5.25e-13
+ AS=5.25e-13 PD=1.021e-05 PS=1.021e-05 M=1 sca=5.3309 scb=0.00475363
+ scc=0.000349818 lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XX289/D0_noxref VSS VDD diodenwx  AREA=6.83795e-12 perim=1.233e-05 sizedup=0
XX289/D1_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D2_noxref VSS VDD diodenwx  AREA=6.83795e-12 perim=1.233e-05 sizedup=0
XX289/D3_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D4_noxref VSS VDD diodenwx  AREA=6.83795e-12 perim=1.233e-05 sizedup=0
XX289/D5_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D6_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D7_noxref VSS VDD diodenwx  AREA=6.83795e-12 perim=1.233e-05 sizedup=0
XX289/D8_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D9_noxref VSS VDD diodenwx  AREA=2.26921e-11 perim=1.915e-05 sizedup=0
XX289/D10_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D11_noxref VSS VDD diodenwx  AREA=2.26921e-11 perim=1.915e-05 sizedup=0
XX289/D12_noxref VSS VDD diodenwx  AREA=6.83795e-12 perim=1.233e-05 sizedup=0
XX289/D13_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D14_noxref VSS VDD diodenwx  AREA=6.83795e-12 perim=1.233e-05 sizedup=0
XX289/D15_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D16_noxref VSS VDD diodenwx  AREA=6.83795e-12 perim=1.233e-05 sizedup=0
XX289/D17_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D18_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D19_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D20_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D21_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D22_noxref VSS VDD diodenwx  AREA=8.8431e-12 perim=1.32e-05 sizedup=0
XX289/D23_noxref VSS VDD diodenwx  AREA=9.97645e-11 perim=4.508e-05 sizedup=0
XX289/D24_noxref VSS VDD diodenwx  AREA=1.69725e-11 perim=1.66e-05 sizedup=0
XXI12/XG1/M2 XI12/N2 DOI VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=1.43975 scb=0.000221266 scc=8.52026e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI12/XG2/M2 XI12/N3 XI12/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.89e-13 PD=3.81e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG3/M2 XI12/N4 XI12/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.89e-13 PD=1.92e-06 PS=3.81e-06 M=1 sca=2.30009 scb=0.000378829
+ scc=4.60368e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG3/M2@3 XI12/N4 XI12/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=2.30009 scb=0.000378829
+ scc=4.60368e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=2.55e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG3/M2@2 XI12/N4 XI12/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.08e-13 PD=3.81e-06 PS=1.92e-06 M=1 sca=2.30009 scb=0.000378829
+ scc=4.60368e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=4.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M2 DLBI XI12/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.89e-13
+ PD=1.92e-06 PS=3.81e-06 M=1 sca=2.30009 scb=0.000378829 scc=4.60368e-07
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07 sb=1.305e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI12/XG4/M2@9 DLBI XI12/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=2.30009 scb=0.000378829
+ scc=4.60368e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=2.55e-07
+ sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M2@8 DLBI XI12/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=2.30009 scb=0.000378829
+ scc=4.60368e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=4.05e-07
+ sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M2@7 DLBI XI12/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=2.30009 scb=0.000378829
+ scc=4.60368e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=5.55e-07
+ sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M2@6 DLBI XI12/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=2.30009 scb=0.000378829
+ scc=4.60368e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=7.05e-07
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M2@5 DLBI XI12/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=2.30009 scb=0.000378829
+ scc=4.60368e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=8.55e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M2@4 DLBI XI12/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=2.30009 scb=0.000378829
+ scc=4.60368e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.005e-06
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M2@3 DLBI XI12/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=2.30009 scb=0.000378829
+ scc=4.60368e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.155e-06
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M2@2 DLBI XI12/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.08e-13 PD=3.81e-06 PS=1.92e-06 M=1 sca=2.30009 scb=0.000378829
+ scc=4.60368e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.305e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI9A0/XG1/M2 XI9A0/N2 CA0 VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=4.07535 scb=0.00152294 scc=2.83909e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI9A0/XG2/M2 CAI0 XI9A0/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.89e-13 PD=3.81e-06 PS=3.81e-06 M=1 sca=2.76719 scb=0.000520562
+ scc=2.85852e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI9A1/XG1/M2 XI9A1/N2 CA1 VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=1.43975 scb=0.000221266 scc=8.52026e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI9A1/XG2/M2 CAI1 XI9A1/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.89e-13 PD=3.81e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI9A2/XG1/M2 XI9A2/N2 CA2 VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=1.43975 scb=0.000221266 scc=8.52026e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI9A2/XG2/M2 CAI2 XI9A2/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.89e-13 PD=3.81e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI8/XG1/M2 XI8/N2 PD VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=1.43975 scb=0.000221266 scc=8.52026e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI8/XG2/M2 PDI XI8/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13 AS=1.89e-13
+ PD=3.81e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05 scc=2.87106e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI6/X1I81/M3 XI6/N0 PDI VSS VSS nfet L=3e-08 W=1.1e-07 AD=6.6e-15 AS=1.265e-14
+ PD=2.3e-07 PS=4.5e-07 M=1 sca=3.70486 scb=0.00288287 scc=1.62404e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9.9e-08 sa=1.15e-07 sb=2.65e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI6/X1I81/M4 XI6/N0 PDTX VSS VSS nfet L=3e-08 W=1.1e-07 AD=6.6e-15 AS=1.265e-14
+ PD=2.3e-07 PS=4.5e-07 M=1 sca=3.70486 scb=0.00288287 scc=1.62404e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9.9e-08 sa=2.65e-07 sb=1.15e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI6/XG0/M2 XI6/N1 XI6/N0 VSS VSS nfet L=3e-08 W=4e-07 AD=4.4e-14 AS=4.4e-14
+ PD=1.02e-06 PS=1.02e-06 M=1 sca=3.05172 scb=0.00191169 scc=7.66588e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.6e-07 sa=1.1e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI6/XG1/M2 XI6/N2 XI6/N1 VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=2.72091 scb=0.00149505 scc=5.33085e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI6/XG2/M2 XI6/N3 XI6/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13 AS=1.89e-13
+ PD=3.81e-06 PS=3.81e-06 M=1 sca=1.64863 scb=0.00056999 scc=1.79823e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI6/XG3/M2 XI6/N4 XI6/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.89e-13
+ PD=1.92e-06 PS=3.81e-06 M=1 sca=1.64863 scb=0.00056999 scc=1.79823e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI6/XG3/M2@3 XI6/N4 XI6/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=2.55e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG3/M2@2 XI6/N4 XI6/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.08e-13 PD=3.81e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=4.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M2 PDTXI XI6/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.89e-13
+ PD=1.92e-06 PS=3.81e-06 M=1 sca=1.64863 scb=0.00056999 scc=1.79823e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07 sb=1.305e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI6/XG4/M2@9 PDTXI XI6/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=2.55e-07
+ sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M2@8 PDTXI XI6/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=4.05e-07
+ sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M2@7 PDTXI XI6/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=5.55e-07
+ sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M2@6 PDTXI XI6/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=7.05e-07
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M2@5 PDTXI XI6/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=8.55e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M2@4 PDTXI XI6/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.005e-06
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M2@3 PDTXI XI6/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.155e-06
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M2@2 PDTXI XI6/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.08e-13 PD=3.81e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.305e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/X1I81/M3 XI7/N0 PDI VSS VSS nfet L=3e-08 W=1.1e-07 AD=6.6e-15 AS=1.265e-14
+ PD=2.3e-07 PS=4.5e-07 M=1 sca=3.70486 scb=0.00288287 scc=1.62404e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9.9e-08 sa=1.15e-07 sb=2.65e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI7/X1I81/M4 XI7/N0 PDRX VSS VSS nfet L=3e-08 W=1.1e-07 AD=6.6e-15 AS=1.265e-14
+ PD=2.3e-07 PS=4.5e-07 M=1 sca=3.70486 scb=0.00288287 scc=1.62404e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9.9e-08 sa=2.65e-07 sb=1.15e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI7/XG0/M2 XI7/N1 XI7/N0 VSS VSS nfet L=3e-08 W=4e-07 AD=4.4e-14 AS=4.4e-14
+ PD=1.02e-06 PS=1.02e-06 M=1 sca=3.05172 scb=0.00191169 scc=7.66588e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.6e-07 sa=1.1e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI7/XG1/M2 XI7/N2 XI7/N1 VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=2.72091 scb=0.00149505 scc=5.33085e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI7/XG2/M2 XI7/N3 XI7/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13 AS=1.89e-13
+ PD=3.81e-06 PS=3.81e-06 M=1 sca=1.64863 scb=0.00056999 scc=1.79823e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI7/XG3/M2 XI7/N4 XI7/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.89e-13
+ PD=1.92e-06 PS=3.81e-06 M=1 sca=1.64863 scb=0.00056999 scc=1.79823e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI7/XG3/M2@3 XI7/N4 XI7/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=2.55e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG3/M2@2 XI7/N4 XI7/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.08e-13 PD=3.81e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=4.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M2 PDRXI XI7/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.89e-13
+ PD=1.92e-06 PS=3.81e-06 M=1 sca=1.64863 scb=0.00056999 scc=1.79823e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07 sb=1.305e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI7/XG4/M2@9 PDRXI XI7/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=2.55e-07
+ sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M2@8 PDRXI XI7/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=4.05e-07
+ sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M2@7 PDRXI XI7/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=5.55e-07
+ sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M2@6 PDRXI XI7/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=7.05e-07
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M2@5 PDRXI XI7/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=8.55e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M2@4 PDRXI XI7/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.005e-06
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M2@3 PDRXI XI7/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.155e-06
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M2@2 PDRXI XI7/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.08e-13 PD=3.81e-06 PS=1.92e-06 M=1 sca=1.64863 scb=0.00056999
+ scc=1.79823e-06 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.305e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG1/M2 XI11/N2 DLBI VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=1.43975 scb=0.000221266 scc=8.52026e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI11/XG2/M2 XI11/N3 XI11/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.89e-13 PD=3.81e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG3/M2 XI11/N4 XI11/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.89e-13 PD=1.92e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG3/M2@3 XI11/N4 XI11/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=2.55e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG3/M2@2 XI11/N4 XI11/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.08e-13 PD=3.81e-06 PS=1.92e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=4.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M2 DLB XI11/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.89e-13
+ PD=1.92e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05 scc=2.87106e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07 sb=1.305e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI11/XG4/M2@9 DLB XI11/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=2.55e-07
+ sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M2@8 DLB XI11/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=4.05e-07
+ sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M2@7 DLB XI11/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=5.55e-07
+ sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M2@6 DLB XI11/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=7.05e-07
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M2@5 DLB XI11/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=8.55e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M2@4 DLB XI11/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.005e-06
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M2@3 DLB XI11/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=2.05471 scb=0.000150854
+ scc=3.34714e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.155e-06
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M2@2 DLB XI11/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.08e-13 PD=3.81e-06 PS=1.92e-06 M=1 sca=2.20617 scb=0.000198572
+ scc=4.35247e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.305e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI5A0/XG1/M2 XI5A0/N2 CCM0 VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=1.43975 scb=0.000221266 scc=8.52026e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI5A0/XG2/M2 CCMI0 XI5A0/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.89e-13 PD=3.81e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI5A1/XG1/M2 XI5A1/N2 CCM1 VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=1.43975 scb=0.000221266 scc=8.52026e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI5A1/XG2/M2 CCMI1 XI5A1/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.89e-13 PD=3.81e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI5A2/XG1/M2 XI5A2/N2 CCM2 VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=1.43975 scb=0.000221266 scc=8.52026e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI5A2/XG2/M2 CCMI2 XI5A2/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.89e-13 PD=3.81e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI3/X1I242/M2 N1N291 XI3/N1 VSS VSS nfet L=3e-08 W=5e-07 AD=5.25e-14
+ AS=5.25e-14 PD=1.21e-06 PS=1.21e-06 M=1 sca=1.50221 scb=0.000250162
+ scc=1.00975e-07 lpccnr=3.1e-08 covpccnr=0 wrxcnr=4.5e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI3/XG0/M3 XI3/N1 DLB XI3/XG0/N1 VSS nfet L=3e-08 W=1e-06 AD=1.1e-13
+ AS=6.75e-14 PD=2.22e-06 PS=1.135e-06 M=1 sca=1.1749 scb=0.000120572
+ scc=3.42144e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=1.1e-07 sb=2.75e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI3/XG0/M4 XI3/XG0/N1 LBEN VSS VSS nfet L=3e-08 W=1e-06 AD=6.75e-14 AS=1.1e-13
+ PD=1.135e-06 PS=2.22e-06 M=1 sca=1.1749 scb=0.000120572 scc=3.42144e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=2.75e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG0A/M2 XI4/SLB LBEN VSS VSS nfet L=3e-08 W=4e-07 AD=4.4e-14 AS=4.4e-14
+ PD=1.02e-06 PS=1.02e-06 M=1 sca=1.48682 scb=0.00023539 scc=8.13879e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.6e-07 sa=1.1e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG0B/M2 XI4/SL XI4/SLB VSS VSS nfet L=3e-08 W=4e-07 AD=4.4e-14 AS=4.4e-14
+ PD=1.02e-06 PS=1.02e-06 M=1 sca=1.48682 scb=0.00023539 scc=8.13879e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.6e-07 sa=1.1e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG0/M4 XI4/XG0/N1 XI4/SLB VSS VSS nfet L=3e-08 W=1e-06 AD=6.75e-14
+ AS=1.1e-13 PD=1.135e-06 PS=2.22e-06 M=1 sca=1.1749 scb=0.000120572
+ scc=3.42144e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=1.1e-07 sb=2.75e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI4/XG0/M3 XI4/N1 DI XI4/XG0/N1 VSS nfet L=3e-08 W=1e-06 AD=1.1e-13 AS=6.75e-14
+ PD=2.22e-06 PS=1.135e-06 M=1 sca=1.1749 scb=0.000120572 scc=3.42144e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=2.75e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG2/M3 DTX XI4/N1 XI4/XG2/N1 VSS nfet L=3e-08 W=2e-06 AD=2.2e-13 AS=1.4e-13
+ PD=4.22e-06 PS=2.14e-06 M=1 sca=0.870522 scb=6.19181e-05 scc=1.71159e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.1e-07 sb=2.8e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG2/M4 XI4/XG2/N1 XI4/N2 VSS VSS nfet L=3e-08 W=2e-06 AD=1.4e-13 AS=2.2e-13
+ PD=2.14e-06 PS=4.22e-06 M=1 sca=0.870522 scb=6.19181e-05 scc=1.71159e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.8e-06 sa=2.8e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG1/M3 XI4/N2 N1N291 XI4/XG1/N1 VSS nfet L=3e-08 W=1e-06 AD=1.1e-13
+ AS=6.75e-14 PD=2.22e-06 PS=1.135e-06 M=1 sca=1.1749 scb=0.000120572
+ scc=3.42144e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=1.1e-07 sb=2.75e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI4/XG1/M4 XI4/XG1/N1 XI4/SL VSS VSS nfet L=3e-08 W=1e-06 AD=6.75e-14
+ AS=1.1e-13 PD=1.135e-06 PS=2.22e-06 M=1 sca=1.1749 scb=0.000120572
+ scc=3.42144e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=2.75e-07 sb=1.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI12/XG1/M1 XI12/N2 DOI VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13 AS=1.26e-13
+ PD=2.61e-06 PS=2.61e-06 M=1 sca=20.544 scb=0.0159143 scc=0.00253599
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI12/XG2/M1 XI12/N3 XI12/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=3.78e-13 PD=7.41e-06 PS=7.41e-06 M=1 sca=9.18389 scb=0.00636638
+ scc=0.000856992 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG3/M1 XI12/N4 XI12/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=3.78e-13 PD=3.72e-06 PS=7.41e-06 M=1 sca=10.3654 scb=0.00645938
+ scc=0.000857001 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG3/M1@3 XI12/N4 XI12/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=10.536 scb=0.00652478
+ scc=0.000857021 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=2.55e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG3/M1@2 XI12/N4 XI12/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=2.16e-13 PD=7.41e-06 PS=3.72e-06 M=1 sca=10.7465 scb=0.00663487
+ scc=0.000857082 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=4.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M1 DLBI XI12/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=3.78e-13
+ PD=3.72e-06 PS=7.41e-06 M=1 sca=11.3985 scb=0.00717751 scc=0.000857972
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07 sb=1.305e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI12/XG4/M1@9 DLBI XI12/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=11.8541 scb=0.00771238
+ scc=0.000859955 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=2.55e-07
+ sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M1@8 DLBI XI12/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=12.4661 scb=0.00857845
+ scc=0.000865867 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=4.05e-07
+ sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M1@7 DLBI XI12/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=13.3156 scb=0.00995883
+ scc=0.000883254 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=5.55e-07
+ sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M1@6 DLBI XI12/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=14.5433 scb=0.0121138
+ scc=0.000933548 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=7.05e-07
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M1@5 DLBI XI12/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=16.412 scb=0.0153839
+ scc=0.00107585 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=8.55e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M1@4 DLBI XI12/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=19.4605 scb=0.0201464
+ scc=0.00146634 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.005e-06
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M1@3 DLBI XI12/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=24.9399 scb=0.0266447
+ scc=0.00249074 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.155e-06
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI12/XG4/M1@2 DLBI XI12/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=2.16e-13 PD=7.41e-06 PS=3.72e-06 M=1 sca=36.3371 scb=0.0345142
+ scc=0.00498851 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.305e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC0@67 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@66 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@65 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@64 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@63 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@62 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@61 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@60 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@59 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI9A0/XG1/M1 XI9A0/N2 CA0 VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13
+ AS=1.26e-13 PD=2.61e-06 PS=2.61e-06 M=1 sca=47.2086 scb=0.0491374
+ scc=0.00508856 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI9A0/XG2/M1 CAI0 XI9A0/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=3.78e-13 PD=7.41e-06 PS=7.41e-06 M=1 sca=36.8462 scb=0.0400538
+ scc=0.00366829 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC0@58 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@57 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI9A1/XG1/M1 XI9A1/N2 CA1 VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13
+ AS=1.26e-13 PD=2.61e-06 PS=2.61e-06 M=1 sca=47.2086 scb=0.0491374
+ scc=0.00508856 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI9A1/XG2/M1 CAI1 XI9A1/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=3.78e-13 PD=7.41e-06 PS=7.41e-06 M=1 sca=36.8462 scb=0.0400538
+ scc=0.00366829 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC0@56 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@55 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI9A2/XG1/M1 XI9A2/N2 CA2 VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13
+ AS=1.26e-13 PD=2.61e-06 PS=2.61e-06 M=1 sca=47.2086 scb=0.0491374
+ scc=0.00508856 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI9A2/XG2/M1 CAI2 XI9A2/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=3.78e-13 PD=7.41e-06 PS=7.41e-06 M=1 sca=36.8462 scb=0.0400538
+ scc=0.00366829 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC0@54 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@53 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@52 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@51 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI8/XG1/M1 XI8/N2 PD VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13 AS=1.26e-13
+ PD=2.61e-06 PS=2.61e-06 M=1 sca=47.2086 scb=0.0491374 scc=0.00508856
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI8/XG2/M1 PDI XI8/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13 AS=3.78e-13
+ PD=7.41e-06 PS=7.41e-06 M=1 sca=36.8462 scb=0.0400538 scc=0.00366829
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI6/X1I81/M1 XI6/X1I81/N1 PDI VDD VDD pfet L=3e-08 W=8e-07 AD=4.8e-14
+ AS=8.4e-14 PD=9.2e-07 PS=1.81e-06 M=1 sca=25.0645 scb=0.0292013 scc=0.00265586
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=7.2e-07 sa=1.05e-07 sb=2.55e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI6/X1I81/M2 XI6/N0 PDTX XI6/X1I81/N1 VDD pfet L=3e-08 W=8e-07 AD=8.4e-14
+ AS=4.8e-14 PD=1.81e-06 PS=9.2e-07 M=1 sca=17.5242 scb=0.0219489 scc=0.00108476
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=7.2e-07 sa=2.55e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI6/XG0/M1 XI6/N1 XI6/N0 VDD VDD pfet L=3e-08 W=8e-07 AD=8.8e-14 AS=8.8e-14
+ PD=1.82e-06 PS=1.82e-06 M=1 sca=10.9 scb=0.0118478 scc=0.000215318
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=7.2e-07 sa=1.1e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC0@50 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@49 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI6/XG1/M1 XI6/N2 XI6/N1 VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13 AS=1.26e-13
+ PD=2.61e-06 PS=2.61e-06 M=1 sca=7.41366 scb=0.00606487 scc=8.56364e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI6/XG2/M1 XI6/N3 XI6/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13 AS=3.78e-13
+ PD=7.41e-06 PS=7.41e-06 M=1 sca=5.59581 scb=0.00296718 scc=3.76795e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI6/XG3/M1 XI6/N4 XI6/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=3.78e-13
+ PD=3.72e-06 PS=7.41e-06 M=1 sca=6.13595 scb=0.00253546 scc=3.68624e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI6/XG3/M1@3 XI6/N4 XI6/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=6.09915 scb=0.00249451
+ scc=3.68256e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=2.55e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG3/M1@2 XI6/N4 XI6/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=2.16e-13 PD=7.41e-06 PS=3.72e-06 M=1 sca=6.14125 scb=0.00254144
+ scc=3.68682e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=4.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M1 PDTXI XI6/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=3.78e-13
+ PD=3.72e-06 PS=7.41e-06 M=1 sca=5.62195 scb=0.00299434 scc=3.77495e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07 sb=1.305e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI6/XG4/M1@9 PDTXI XI6/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=6.07751 scb=0.00352921
+ scc=3.97331e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=2.55e-07
+ sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M1@8 PDTXI XI6/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=6.6896 scb=0.00439528
+ scc=4.56445e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=4.05e-07
+ sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M1@7 PDTXI XI6/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=7.5391 scb=0.00577566
+ scc=6.30318e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=5.55e-07
+ sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M1@6 PDTXI XI6/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=8.76674 scb=0.00793061
+ scc=0.000113325 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=7.05e-07
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M1@5 PDTXI XI6/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=10.6355 scb=0.0112007
+ scc=0.000255623 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=8.55e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M1@4 PDTXI XI6/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=13.684 scb=0.0159632
+ scc=0.000646117 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.005e-06
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M1@3 PDTXI XI6/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=19.1633 scb=0.0224615
+ scc=0.00167052 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.155e-06
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI6/XG4/M1@2 PDTXI XI6/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=2.16e-13 PD=7.41e-06 PS=3.72e-06 M=1 sca=30.5606 scb=0.030331
+ scc=0.00416829 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.305e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC0@48 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@47 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI7/X1I81/M1 XI7/X1I81/N1 PDI VDD VDD pfet L=3e-08 W=8e-07 AD=4.8e-14
+ AS=8.4e-14 PD=9.2e-07 PS=1.81e-06 M=1 sca=25.0645 scb=0.0292013 scc=0.00265586
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=7.2e-07 sa=1.05e-07 sb=2.55e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI7/X1I81/M2 XI7/N0 PDRX XI7/X1I81/N1 VDD pfet L=3e-08 W=8e-07 AD=8.4e-14
+ AS=4.8e-14 PD=1.81e-06 PS=9.2e-07 M=1 sca=17.5242 scb=0.0219489 scc=0.00108476
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=7.2e-07 sa=2.55e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI7/XG0/M1 XI7/N1 XI7/N0 VDD VDD pfet L=3e-08 W=8e-07 AD=8.8e-14 AS=8.8e-14
+ PD=1.82e-06 PS=1.82e-06 M=1 sca=10.9 scb=0.0118478 scc=0.000215318
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=7.2e-07 sa=1.1e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI7/XG1/M1 XI7/N2 XI7/N1 VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13 AS=1.26e-13
+ PD=2.61e-06 PS=2.61e-06 M=1 sca=7.41366 scb=0.00606487 scc=8.56364e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI7/XG2/M1 XI7/N3 XI7/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13 AS=3.78e-13
+ PD=7.41e-06 PS=7.41e-06 M=1 sca=5.59581 scb=0.00296718 scc=3.76795e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI7/XG3/M1 XI7/N4 XI7/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=3.78e-13
+ PD=3.72e-06 PS=7.41e-06 M=1 sca=6.13595 scb=0.00253546 scc=3.68624e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI7/XG3/M1@3 XI7/N4 XI7/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=6.09915 scb=0.00249451
+ scc=3.68256e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=2.55e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG3/M1@2 XI7/N4 XI7/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=2.16e-13 PD=7.41e-06 PS=3.72e-06 M=1 sca=6.14125 scb=0.00254144
+ scc=3.68682e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=4.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M1 PDRXI XI7/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=3.78e-13
+ PD=3.72e-06 PS=7.41e-06 M=1 sca=5.62195 scb=0.00299434 scc=3.77495e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07 sb=1.305e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI7/XG4/M1@9 PDRXI XI7/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=6.07751 scb=0.00352921
+ scc=3.97331e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=2.55e-07
+ sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M1@8 PDRXI XI7/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=6.6896 scb=0.00439528
+ scc=4.56445e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=4.05e-07
+ sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M1@7 PDRXI XI7/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=7.5391 scb=0.00577566
+ scc=6.30318e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=5.55e-07
+ sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M1@6 PDRXI XI7/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=8.76674 scb=0.00793061
+ scc=0.000113325 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=7.05e-07
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M1@5 PDRXI XI7/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=10.6355 scb=0.0112007
+ scc=0.000255623 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=8.55e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M1@4 PDRXI XI7/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=13.684 scb=0.0159632
+ scc=0.000646117 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.005e-06
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M1@3 PDRXI XI7/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=19.1633 scb=0.0224615
+ scc=0.00167052 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.155e-06
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI7/XG4/M1@2 PDRXI XI7/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=2.16e-13 PD=7.41e-06 PS=3.72e-06 M=1 sca=30.5606 scb=0.030331
+ scc=0.00416829 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.305e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG1/M1 XI11/N2 DLBI VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13 AS=1.26e-13
+ PD=2.61e-06 PS=2.61e-06 M=1 sca=40.4882 scb=0.0397626 scc=0.00507805
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI11/XG2/M1 XI11/N3 XI11/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=3.78e-13 PD=7.41e-06 PS=7.41e-06 M=1 sca=17.257 scb=0.0167881
+ scc=0.00116592 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG3/M1 XI11/N4 XI11/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=3.78e-13 PD=3.72e-06 PS=7.41e-06 M=1 sca=14.7064 scb=0.010411
+ scc=0.000889573 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG3/M1@3 XI11/N4 XI11/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=13.9658 scb=0.00896466
+ scc=0.000868058 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=2.55e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG3/M1@2 XI11/N4 XI11/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=2.16e-13 PD=7.41e-06 PS=3.72e-06 M=1 sca=13.5245 scb=0.00812271
+ scc=0.000860776 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=4.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M1 DLB XI11/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=3.78e-13
+ PD=3.72e-06 PS=7.41e-06 M=1 sca=13.2855 scb=0.00767946 scc=0.000858318
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07 sb=1.305e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI11/XG4/M1@9 DLB XI11/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=13.4646 scb=0.00801056
+ scc=0.000860068 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=2.55e-07
+ sb=1.155e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M1@8 DLB XI11/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=13.8568 scb=0.00875456
+ scc=0.000865903 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=4.05e-07
+ sb=1.005e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M1@7 DLB XI11/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=14.5286 scb=0.0100623
+ scc=0.000883266 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=5.55e-07
+ sb=8.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M1@6 DLB XI11/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=15.6105 scb=0.0121743
+ scc=0.000933551 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=7.05e-07
+ sb=7.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M1@5 DLB XI11/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=16.412 scb=0.0153839
+ scc=0.00107585 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=8.55e-07
+ sb=5.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M1@4 DLB XI11/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=19.4605 scb=0.0201464
+ scc=0.00146634 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.005e-06
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M1@3 DLB XI11/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=24.9399 scb=0.0266447
+ scc=0.00249074 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.155e-06
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI11/XG4/M1@2 DLB XI11/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=2.16e-13 PD=7.41e-06 PS=3.72e-06 M=1 sca=36.3371 scb=0.0345142
+ scc=0.00498851 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.305e-06
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC0@46 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@45 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@44 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@43 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@42 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@41 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@40 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@39 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@38 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@37 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@36 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@35 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@34 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@33 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@32 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI5A0/XG1/M1 XI5A0/N2 CCM0 VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13
+ AS=1.26e-13 PD=2.61e-06 PS=2.61e-06 M=1 sca=47.2086 scb=0.0491374
+ scc=0.00508856 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI5A0/XG2/M1 CCMI0 XI5A0/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=3.78e-13 PD=7.41e-06 PS=7.41e-06 M=1 sca=36.8462 scb=0.0400538
+ scc=0.00366829 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC0@31 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@30 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI5A1/XG1/M1 XI5A1/N2 CCM1 VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13
+ AS=1.26e-13 PD=2.61e-06 PS=2.61e-06 M=1 sca=47.2086 scb=0.0491374
+ scc=0.00508856 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI5A1/XG2/M1 CCMI1 XI5A1/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=3.78e-13 PD=7.41e-06 PS=7.41e-06 M=1 sca=36.8462 scb=0.0400538
+ scc=0.00366829 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC0@29 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@28 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI5A2/XG1/M1 XI5A2/N2 CCM2 VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13
+ AS=1.26e-13 PD=2.61e-06 PS=2.61e-06 M=1 sca=47.2086 scb=0.0491374
+ scc=0.00508856 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI5A2/XG2/M1 CCMI2 XI5A2/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=3.78e-13 PD=7.41e-06 PS=7.41e-06 M=1 sca=36.8462 scb=0.0400538
+ scc=0.00366829 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XMDC0@27 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@26 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@25 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@24 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@23 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@22 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@21 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@20 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@19 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@18 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI3/X1I242/M1 N1N291 XI3/N1 VDD VDD pfet L=3e-08 W=1e-06 AD=1.05e-13
+ AS=1.05e-13 PD=2.21e-06 PS=2.21e-06 M=1 sca=40.515 scb=0.0389876 scc=0.003988
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI3/XG0/M1 XI3/N1 DLB VDD VDD pfet L=3e-08 W=1e-06 AD=6.75e-14 AS=1.1e-13
+ PD=1.135e-06 PS=2.22e-06 M=1 sca=48.1006 scb=0.0380682 scc=0.00444314
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=1.1e-07 sb=2.75e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI3/XG0/M2 XI3/N1 LBEN VDD VDD pfet L=3e-08 W=1e-06 AD=6.75e-14 AS=1.1e-13
+ PD=1.135e-06 PS=2.22e-06 M=1 sca=51.432 scb=0.0419461 scc=0.00516742
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=2.75e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC0@17 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@16 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=7.41019 scb=0.00658528 scc=0.000443878
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI4/XG0A/M1 XI4/SLB LBEN VDD VDD pfet L=3e-08 W=8e-07 AD=8.8e-14 AS=8.8e-14
+ PD=1.82e-06 PS=1.82e-06 M=1 sca=51.3739 scb=0.0381234 scc=0.00559503
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=7.2e-07 sa=1.1e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG0B/M1 XI4/SL XI4/SLB VDD VDD pfet L=3e-08 W=8e-07 AD=8.8e-14 AS=8.8e-14
+ PD=1.82e-06 PS=1.82e-06 M=1 sca=45.8097 scb=0.0290937 scc=0.00498534
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=7.2e-07 sa=1.1e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG0/M2 XI4/N1 XI4/SLB VDD VDD pfet L=3e-08 W=1e-06 AD=6.75e-14 AS=1.1e-13
+ PD=1.135e-06 PS=2.22e-06 M=1 sca=37.9537 scb=0.0221736 scc=0.00396158
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=1.1e-07 sb=2.75e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG0/M1 XI4/N1 DI VDD VDD pfet L=3e-08 W=1e-06 AD=6.75e-14 AS=1.1e-13
+ PD=1.135e-06 PS=2.22e-06 M=1 sca=37.5879 scb=0.0215191 scc=0.00395775
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=2.75e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG2/M1 DTX XI4/N1 VDD VDD pfet L=3e-08 W=2e-06 AD=1.4e-13 AS=2.2e-13
+ PD=2.14e-06 PS=4.22e-06 M=1 sca=23.1954 scb=0.0132161 scc=0.00199092
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.8e-06 sa=1.1e-07 sb=2.8e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG2/M2 DTX XI4/N2 VDD VDD pfet L=3e-08 W=2e-06 AD=1.4e-13 AS=2.2e-13
+ PD=2.14e-06 PS=4.22e-06 M=1 sca=24.0579 scb=0.0148627 scc=0.00201478
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.8e-06 sa=2.8e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG1/M1 XI4/N2 N1N291 VDD VDD pfet L=3e-08 W=1e-06 AD=6.75e-14 AS=1.1e-13
+ PD=1.135e-06 PS=2.22e-06 M=1 sca=42.2268 scb=0.0314477 scc=0.00432264
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=1.1e-07 sb=2.75e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI4/XG1/M2 XI4/N2 XI4/SL VDD VDD pfet L=3e-08 W=1e-06 AD=6.75e-14 AS=1.1e-13
+ PD=1.135e-06 PS=2.22e-06 M=1 sca=46.8083 scb=0.0377287 scc=0.00506335
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=9e-07 sa=2.75e-07 sb=1.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XMDC0@15 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@14 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@13 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@12 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@11 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@10 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@9 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@8 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@7 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@6 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@5 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@4 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@3 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XMDC0@2 VDD VSS VDD VDD pfet L=5e-06 W=5e-06 AD=5.25e-13 AS=5.25e-13
+ PD=1.021e-05 PS=1.021e-05 M=1 sca=4.30942 scb=0.00379615 scc=0.000194942
+ lpccnr=4.504e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG1/M2 XI10/N2 DOI VSS VSS nfet L=3e-08 W=6e-07 AD=6.3e-14 AS=6.3e-14
+ PD=1.41e-06 PS=1.41e-06 M=1 sca=1.43975 scb=0.000221266 scc=8.52026e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.4e-07 sa=1.05e-07 sb=1.05e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI10/XG2/M2 XI10/N3 XI10/N2 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.89e-13 PD=3.81e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI10/XG3/M2 XI10/N4 XI10/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.89e-13 PD=1.92e-06 PS=3.81e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI10/XG3/M2@3 XI10/N4 XI10/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13
+ AS=1.08e-13 PD=1.92e-06 PS=1.92e-06 M=1 sca=0.9605 scb=8.34304e-05
+ scc=2.87106e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=2.55e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI10/XG3/M2@2 XI10/N4 XI10/N3 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13
+ AS=1.08e-13 PD=3.81e-06 PS=1.92e-06 M=1 sca=1.52348 scb=0.000117647
+ scc=3.10788e-08 lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=4.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI10/XG4/M2 DO XI10/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.89e-13
+ PD=1.92e-06 PS=3.81e-06 M=1 sca=1.71053 scb=0.000190051 scc=5.52515e-08
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.05e-07 sb=1.305e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M2@9 DO XI10/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.08e-13
+ PD=1.92e-06 PS=1.92e-06 M=1 sca=1.83198 scb=0.00026366 scc=1.10458e-07
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=2.55e-07 sb=1.155e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M2@8 DO XI10/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.08e-13
+ PD=1.92e-06 PS=1.92e-06 M=1 sca=1.9855 scb=0.000386237 scc=2.78965e-07
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=4.05e-07 sb=1.005e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M2@7 DO XI10/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.08e-13
+ PD=1.92e-06 PS=1.92e-06 M=1 sca=2.18348 scb=0.000588545 scc=7.89347e-07
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=5.55e-07 sb=8.55e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M2@6 DO XI10/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.08e-13
+ PD=1.92e-06 PS=1.92e-06 M=1 sca=2.4449 scb=0.000918836 scc=2.32091e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=7.05e-07 sb=7.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M2@5 DO XI10/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.08e-13
+ PD=1.92e-06 PS=1.92e-06 M=1 sca=2.80006 scb=0.00145081 scc=6.86484e-06
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=8.55e-07 sb=5.55e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M2@4 DO XI10/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.08e-13
+ PD=1.92e-06 PS=1.92e-06 M=1 sca=3.2998 scb=0.00229283 scc=2.01548e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.005e-06 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M2@3 DO XI10/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.08e-13 AS=1.08e-13
+ PD=1.92e-06 PS=1.92e-06 M=1 sca=4.03473 scb=0.00359515 scc=5.83151e-05
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.155e-06 sb=2.55e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M2@2 DO XI10/N4 VSS VSS nfet L=3e-08 W=1.8e-06 AD=1.89e-13 AS=1.08e-13
+ PD=3.81e-06 PS=1.92e-06 M=1 sca=5.17943 scb=0.00554553 scc=0.00016521
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.62e-06 sa=1.305e-06 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG1/M1 XI10/N2 DOI VDD VDD pfet L=3e-08 W=1.2e-06 AD=1.26e-13 AS=1.26e-13
+ PD=2.61e-06 PS=2.61e-06 M=1 sca=20.544 scb=0.0159143 scc=0.00253599
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=1.08e-06 sa=1.05e-07 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG2/M1 XI10/N3 XI10/N2 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=3.78e-13 PD=7.41e-06 PS=7.41e-06 M=1 sca=9.18389 scb=0.00636638
+ scc=0.000856992 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI10/XG3/M1 XI10/N4 XI10/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=3.78e-13 PD=3.72e-06 PS=7.41e-06 M=1 sca=10.3654 scb=0.00645938
+ scc=0.000857001 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07
+ sb=4.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI10/XG3/M1@3 XI10/N4 XI10/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13
+ AS=2.16e-13 PD=3.72e-06 PS=3.72e-06 M=1 sca=10.536 scb=0.00652478
+ scc=0.000857021 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=2.55e-07
+ sb=2.55e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI10/XG3/M1@2 XI10/N4 XI10/N3 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13
+ AS=2.16e-13 PD=7.41e-06 PS=3.72e-06 M=1 sca=10.7465 scb=0.00663487
+ scc=0.000857082 lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=4.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI10/XG4/M1 DO XI10/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=3.78e-13
+ PD=3.72e-06 PS=7.41e-06 M=1 sca=11.3985 scb=0.00717751 scc=0.000857972
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.05e-07 sb=1.305e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M1@9 DO XI10/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=2.16e-13
+ PD=3.72e-06 PS=3.72e-06 M=1 sca=11.8541 scb=0.00771238 scc=0.000859955
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=2.55e-07 sb=1.155e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M1@8 DO XI10/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=2.16e-13
+ PD=3.72e-06 PS=3.72e-06 M=1 sca=12.4661 scb=0.00857845 scc=0.000865867
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=4.05e-07 sb=1.005e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M1@7 DO XI10/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=2.16e-13
+ PD=3.72e-06 PS=3.72e-06 M=1 sca=13.3156 scb=0.00995883 scc=0.000883254
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=5.55e-07 sb=8.55e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M1@6 DO XI10/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=2.16e-13
+ PD=3.72e-06 PS=3.72e-06 M=1 sca=14.5433 scb=0.0121138 scc=0.000933548
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=7.05e-07 sb=7.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M1@5 DO XI10/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=2.16e-13
+ PD=3.72e-06 PS=3.72e-06 M=1 sca=16.412 scb=0.0153839 scc=0.00107585
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=8.55e-07 sb=5.55e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M1@4 DO XI10/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=2.16e-13
+ PD=3.72e-06 PS=3.72e-06 M=1 sca=19.4605 scb=0.0201464 scc=0.00146634
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.005e-06 sb=4.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M1@3 DO XI10/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=2.16e-13 AS=2.16e-13
+ PD=3.72e-06 PS=3.72e-06 M=1 sca=24.9399 scb=0.0266447 scc=0.00249074
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.155e-06 sb=2.55e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI10/XG4/M1@2 DO XI10/N4 VDD VDD pfet L=3e-08 W=3.6e-06 AD=3.78e-13 AS=2.16e-13
+ PD=7.41e-06 PS=3.72e-06 M=1 sca=36.3371 scb=0.0345142 scc=0.00498851
+ lpccnr=3.1e-08 covpccnr=0 wrxcnr=3.24e-06 sa=1.305e-06 sb=1.05e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX290/D0_noxref VSS VDDHA_RX diodenwx  AREA=3.92273e-10 perim=0.00012743
+ sizedup=0
XX290/D1_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782
+ sizedup=0
XX290/D2_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782
+ sizedup=0
XX290/D3_noxref VSS VDDHA_RX diodenwx  AREA=3.3442e-10 perim=0.00012782
+ sizedup=0
XXI2/XI3/M4N XI2/XI3/N3 PDRXI VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=0.960294 scb=3.88199e-05
+ scc=1.62723e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI3/M3N XI2/XI3/N3 PDRXI VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=16.0067 scb=0.0197187
+ scc=0.000873628 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI3/XG2/M1 XI2/PDRXI XI2/XI3/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/XG2/M1@4 XI2/PDRXI XI2/XI3/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/XG2/M1@3 XI2/PDRXI XI2/XI3/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/XG2/M1@2 XI2/PDRXI XI2/XI3/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/XG1/M1 XI2/XI3/N1N36 XI2/XI3/N1N5 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=3.36e-13 AS=3.36e-13 PD=5.84e-06 PS=5.84e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/M3P XI2/XI3/N1N5 XI2/XI3/N2 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=3.43331
+ scb=0.00285132 scc=4.77845e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/M1P XI2/XI3/N2 XI2/XI3/N1 VDDHA_RX VDDHA_RX egpfet L=3e-06 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979 scb=0.00151603
+ scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI3/M1N XI2/XI3/N1 XI2/XI3/N2 VDDHA_RX VDDHA_RX egpfet L=3e-06 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=4.11762 scb=0.0021369
+ scc=3.00661e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI3/XG2/M2 XI2/PDRXI XI2/XI3/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/XG2/M2@4 XI2/PDRXI XI2/XI3/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/XG2/M2@3 XI2/PDRXI XI2/XI3/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/XG2/M2@2 XI2/PDRXI XI2/XI3/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/XG1/M2 XI2/XI3/N1N36 XI2/XI3/N1N5 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/M4P XI2/XI3/N1N5 XI2/XI3/N2 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/M2P XI2/XI3/N2 PDRXI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI3/M2N XI2/XI3/N1 XI2/XI3/N3 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/M4N XI2/XI4/N3 PDTXI VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=0.960294 scb=3.88199e-05
+ scc=1.62723e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI4/M3N XI2/XI4/N3 PDTXI VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=4.43262 scb=0.00417318
+ scc=5.06595e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI4/XG2/M1 XI2/PDTXI XI2/XI4/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/XG2/M1@4 XI2/PDTXI XI2/XI4/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/XG2/M1@3 XI2/PDTXI XI2/XI4/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/XG2/M1@2 XI2/PDTXI XI2/XI4/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/XG1/M1 XI2/XI4/N1N36 XI2/XI4/N1N5 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=3.36e-13 AS=3.36e-13 PD=5.84e-06 PS=5.84e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/M3P XI2/XI4/N1N5 XI2/XI4/N2 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=3.43331
+ scb=0.00285132 scc=4.77845e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/M1P XI2/XI4/N2 XI2/XI4/N1 VDDHA_RX VDDHA_RX egpfet L=3e-06 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979 scb=0.00151603
+ scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI4/M1N XI2/XI4/N1 XI2/XI4/N2 VDDHA_RX VDDHA_RX egpfet L=3e-06 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979 scb=0.00151603
+ scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI4/XG2/M2 XI2/PDTXI XI2/XI4/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/XG2/M2@4 XI2/PDTXI XI2/XI4/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/XG2/M2@3 XI2/PDTXI XI2/XI4/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/XG2/M2@2 XI2/PDTXI XI2/XI4/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/XG1/M2 XI2/XI4/N1N36 XI2/XI4/N1N5 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/M4P XI2/XI4/N1N5 XI2/XI4/N2 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/M2P XI2/XI4/N2 PDTXI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI4/M2N XI2/XI4/N1 XI2/XI4/N3 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/M4N XI2/XI2/N3 PDI VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=0.960294 scb=3.88199e-05
+ scc=1.62723e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI2/M3N XI2/XI2/N3 PDI VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=4.43262 scb=0.00417318
+ scc=5.06595e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI2/XG2/M1 XI2/PDI XI2/XI2/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/XG2/M1@4 XI2/PDI XI2/XI2/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/XG2/M1@3 XI2/PDI XI2/XI2/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/XG2/M1@2 XI2/PDI XI2/XI2/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/XG1/M1 XI2/XI2/N1N36 XI2/XI2/N1N5 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=3.36e-13 AS=3.36e-13 PD=5.84e-06 PS=5.84e-06 M=1 sca=3.39213
+ scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/M3P XI2/XI2/N1N5 XI2/XI2/N2 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=3.43331
+ scb=0.00285132 scc=4.77845e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/M1P XI2/XI2/N2 XI2/XI2/N1 VDDHA_RX VDDHA_RX egpfet L=3e-06 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979 scb=0.00151603
+ scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI2/M1N XI2/XI2/N1 XI2/XI2/N2 VDDHA_RX VDDHA_RX egpfet L=3e-06 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979 scb=0.00151603
+ scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI2/XG2/M2 XI2/PDI XI2/XI2/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/XG2/M2@4 XI2/PDI XI2/XI2/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/XG2/M2@3 XI2/PDI XI2/XI2/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/XG2/M2@2 XI2/PDI XI2/XI2/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/XG1/M2 XI2/XI2/N1N36 XI2/XI2/N1N5 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/M4P XI2/XI2/N1N5 XI2/XI2/N2 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/M2P XI2/XI2/N2 PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI2/M2N XI2/XI2/N1 XI2/XI2/N3 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/M4N XI2/XI5A2/N3 CAI2 VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=0.960294 scb=3.88199e-05
+ scc=1.62723e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI5A2/M3N XI2/XI5A2/N3 CAI2 VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=4.43262 scb=0.00417318
+ scc=5.06595e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI5A2/XG2/M1 XI2/CAI2 XI2/XI5A2/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/XG2/M1@4 XI2/CAI2 XI2/XI5A2/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/XG2/M1@3 XI2/CAI2 XI2/XI5A2/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/XG2/M1@2 XI2/CAI2 XI2/XI5A2/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/XG1/M1 XI2/XI5A2/N1N36 XI2/XI5A2/N1N5 VDDHA_RX VDDHA_RX egpfet
+ L=1.5e-07 W=2.8e-06 AD=3.36e-13 AS=3.36e-13 PD=5.84e-06 PS=5.84e-06 M=1
+ sca=3.39213 scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.52e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/M3P XI2/XI5A2/N1N5 XI2/XI5A2/N2 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=3.43331
+ scb=0.00285132 scc=4.77845e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/M1P XI2/XI5A2/N2 XI2/XI5A2/N1 VDDHA_RX VDDHA_RX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979
+ scb=0.00151603 scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/M1N XI2/XI5A2/N1 XI2/XI5A2/N2 VDDHA_RX VDDHA_RX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979
+ scb=0.00151603 scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/XG2/M2 XI2/CAI2 XI2/XI5A2/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/XG2/M2@4 XI2/CAI2 XI2/XI5A2/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/XG2/M2@3 XI2/CAI2 XI2/XI5A2/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/XG2/M2@2 XI2/CAI2 XI2/XI5A2/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/XG1/M2 XI2/XI5A2/N1N36 XI2/XI5A2/N1N5 VSSA_RX VSSA_RX egnfet
+ L=1.5e-07 W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI5A2/M4P XI2/XI5A2/N1N5 XI2/XI5A2/N2 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/M2P XI2/XI5A2/N2 CAI2 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A2/M2N XI2/XI5A2/N1 XI2/XI5A2/N3 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=6.4e-07 AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI5A1/M4N XI2/XI5A1/N3 CAI1 VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=0.960294 scb=3.88199e-05
+ scc=1.62723e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI5A1/M3N XI2/XI5A1/N3 CAI1 VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=4.43262 scb=0.00417318
+ scc=5.06595e-05 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI5A1/XG2/M1 XI2/CAI1 XI2/XI5A1/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/XG2/M1@4 XI2/CAI1 XI2/XI5A1/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/XG2/M1@3 XI2/CAI1 XI2/XI5A1/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/XG2/M1@2 XI2/CAI1 XI2/XI5A1/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=3.50292
+ scb=0.00329833 scc=0.000163146 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/XG1/M1 XI2/XI5A1/N1N36 XI2/XI5A1/N1N5 VDDHA_RX VDDHA_RX egpfet
+ L=1.5e-07 W=2.8e-06 AD=3.36e-13 AS=3.36e-13 PD=5.84e-06 PS=5.84e-06 M=1
+ sca=3.39213 scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.52e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/M3P XI2/XI5A1/N1N5 XI2/XI5A1/N2 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=3.43331
+ scb=0.00285132 scc=4.77845e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/M1P XI2/XI5A1/N2 XI2/XI5A1/N1 VDDHA_RX VDDHA_RX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979
+ scb=0.00151603 scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/M1N XI2/XI5A1/N1 XI2/XI5A1/N2 VDDHA_RX VDDHA_RX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979
+ scb=0.00151603 scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/XG2/M2 XI2/CAI1 XI2/XI5A1/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/XG2/M2@4 XI2/CAI1 XI2/XI5A1/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/XG2/M2@3 XI2/CAI1 XI2/XI5A1/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/XG2/M2@2 XI2/CAI1 XI2/XI5A1/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/XG1/M2 XI2/XI5A1/N1N36 XI2/XI5A1/N1N5 VSSA_RX VSSA_RX egnfet
+ L=1.5e-07 W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI5A1/M4P XI2/XI5A1/N1N5 XI2/XI5A1/N2 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/M2P XI2/XI5A1/N2 CAI1 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A1/M2N XI2/XI5A1/N1 XI2/XI5A1/N3 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=6.4e-07 AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI5A0/M4N XI2/XI5A0/N3 CAI0 VSS VSS nfet L=3e-08 W=2.8e-07 AD=2.94e-14
+ AS=2.94e-14 PD=7.7e-07 PS=7.7e-07 M=1 sca=0.960294 scb=3.88199e-05
+ scc=1.62723e-09 lpccnr=3.1e-08 covpccnr=0 wrxcnr=2.52e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI5A0/M3N XI2/XI5A0/N3 CAI0 VDD VDD pfet L=3e-08 W=5.6e-07 AD=5.88e-14
+ AS=5.88e-14 PD=1.33e-06 PS=1.33e-06 M=1 sca=12.8857 scb=0.0152062
+ scc=0.000404943 lpccnr=3.1e-08 covpccnr=0 wrxcnr=5.04e-07 sa=1.05e-07
+ sb=1.05e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI5A0/XG2/M1 XI2/CAI0 XI2/XI5A0/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=9.42555
+ scb=0.0100427 scc=0.000276867 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/XG2/M1@4 XI2/CAI0 XI2/XI5A0/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=7.10155
+ scb=0.00601223 scc=0.000177513 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=4.1e-07 sb=7e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/XG2/M1@3 XI2/CAI0 XI2/XI5A0/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=1.96e-13 PD=2.94e-06 PS=2.94e-06 M=1 sca=5.91934
+ scb=0.00433708 scc=0.000164871 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=7e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/XG2/M1@2 XI2/CAI0 XI2/XI5A0/N1N36 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=2.8e-06 AD=1.96e-13 AS=3.36e-13 PD=2.94e-06 PS=5.84e-06 M=1 sca=5.23693
+ scb=0.00368289 scc=0.000163346 lpccnr=1.5e-07 covpccnr=0 wrxcnr=2.52e-06
+ sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/XG1/M1 XI2/XI5A0/N1N36 XI2/XI5A0/N1N5 VDDHA_RX VDDHA_RX egpfet
+ L=1.5e-07 W=2.8e-06 AD=3.36e-13 AS=3.36e-13 PD=5.84e-06 PS=5.84e-06 M=1
+ sca=3.39213 scb=0.00316561 scc=0.000147986 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=2.52e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/M3P XI2/XI5A0/N1N5 XI2/XI5A0/N2 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=3.43331
+ scb=0.00285132 scc=4.77845e-05 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/M1P XI2/XI5A0/N2 XI2/XI5A0/N1 VDDHA_RX VDDHA_RX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979
+ scb=0.00151603 scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/M1N XI2/XI5A0/N1 XI2/XI5A0/N2 VDDHA_RX VDDHA_RX egpfet L=3e-06
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.11979
+ scb=0.00151603 scc=2.94103e-05 lpccnr=2.715e-06 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=2 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/XG2/M2 XI2/CAI0 XI2/XI5A0/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=9.9e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/XG2/M2@4 XI2/CAI0 XI2/XI5A0/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=7e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/XG2/M2@3 XI2/CAI0 XI2/XI5A0/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=5.6e-14 PD=9.4e-07 PS=9.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=7e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/XG2/M2@2 XI2/CAI0 XI2/XI5A0/N1N36 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=8e-07 AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=9.9e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/XG1/M2 XI2/XI5A0/N1N36 XI2/XI5A0/N1N5 VSSA_RX VSSA_RX egnfet
+ L=1.5e-07 W=8e-07 AD=9.6e-14 AS=9.6e-14 PD=1.84e-06 PS=1.84e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI5A0/M4P XI2/XI5A0/N1N5 XI2/XI5A0/N2 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/M2P XI2/XI5A0/N2 CAI0 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=6.4e-07
+ AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI5A0/M2N XI2/XI5A0/N1 XI2/XI5A0/N3 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=6.4e-07 AD=7.68e-14 AS=7.68e-14 PD=1.52e-06 PS=1.52e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=5.76e-07 sa=1.2e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/MDC1@16 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@17 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@18 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@19 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@20 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@21 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@22 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@23 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@24 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@25 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@26 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@27 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@28 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@29 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@30 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@31 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@32 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@33 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@34 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@35 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@36 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@37 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@38 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@39 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@40 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@41 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@42 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@43 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@44 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@45 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@46 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@47 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@48 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@49 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@50 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@51 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@52 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@53 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@54 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@55 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@56 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@57 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@58 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@59 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/MDC1@60 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@2 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@3 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@4 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@5 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@6 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@7 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@8 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@9 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@10 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@11 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@12 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@13 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@14 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@15 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@16 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@17 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@18 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@19 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@20 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@21 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@22 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@23 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@24 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@25 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@26 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@27 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@28 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@29 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@30 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@31 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@32 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@33 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@34 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@35 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@36 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@37 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@38 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@39 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@40 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@41 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@42 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@43 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@44 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@45 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@46 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@47 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@48 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@49 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@50 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@51 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@52 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@53 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@54 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@55 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@56 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@57 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@58 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@59 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/MDCAP2@60 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@2 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@3 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@4 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@5 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@6 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@7 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@8 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@9 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@10 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@11 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@12 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@13 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@14 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@15 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@16 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@17 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@18 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@19 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@20 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@21 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@22 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@23 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@24 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XX290/X12/D0_noxref VSS VDDHA_RX diodenwx  AREA=4.98294e-10 perim=9.888e-05
+ sizedup=0
XXI2/XI1/MDCAP2@25 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.51773 scb=0.00192174
+ scc=9.74806e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@26 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@27 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@28 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=5.25548 scb=0.0046872
+ scc=0.000346407 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@29 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@30 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@31 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@32 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@33 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@34 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@35 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@36 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@37 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@38 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@39 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@40 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@41 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=8.35626 scb=0.00747633
+ scc=0.000595342 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@42 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@43 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@44 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@45 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@46 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@47 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@48 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@49 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@50 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@51 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@52 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@53 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@54 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@55 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/M3 XI2/VBP XI2/XI0/PDB VDDHA_RX VDDHA_RX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=38.4615 scb=0.0292734
+ scc=0.00580942 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/M3@2 XI2/VBP XI2/XI0/PDB VDDHA_RX VDDHA_RX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=6.2475 scb=0.00727366
+ scc=0.000157548 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/MDCAP2@56 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/M1 XI2/N1N12 XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.728e-13 PD=1.58e-06 PS=3.12e-06 M=1 sca=10.3272
+ scb=0.0104019 scc=0.00106356 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06
+ sa=1.2e-07 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/M1@2 XI2/N1N12 XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.728e-13 PD=1.58e-06 PS=3.12e-06 M=1 sca=10.3272
+ scb=0.0104019 scc=0.00106356 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06
+ sa=5.6e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@57 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@58 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/MDCAP2@59 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06
+ AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@2 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/M4 XI2/XI0/INN XI2/XI0/N3 VDDHA_RX VDDHA_RX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.09221 scb=0.000690888
+ scc=7.10442e-07 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/M11 XI2/XI0/PDB XI2/PDI VDDHA_RX VDDHA_RX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=46.6852 scb=0.0399103
+ scc=0.00614241 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI1/MDC1@3 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=6.20155 scb=0.00557825
+ scc=0.000497871 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M27 VDDHA_RX XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=5e-06
+ W=5e-06 AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.35291
+ scb=0.001911 scc=9.74764e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M27@4 VDDHA_RX XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=5e-06
+ W=5e-06 AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471
+ scb=0.00189807 scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M27@3 VDDHA_RX XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=5e-06
+ W=5e-06 AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471
+ scb=0.00189807 scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M27@2 VDDHA_RX XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=5e-06
+ W=5e-06 AD=6e-13 AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=5.25548
+ scb=0.0046872 scc=0.000346407 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M13 XI2/XI0/PDB XI2/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M1 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.728e-13 PD=1.58e-06 PS=3.12e-06 M=1 sca=14.7929
+ scb=0.0126174 scc=0.00176209 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06
+ sa=1.2e-07 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M2 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.728e-13 PD=1.58e-06 PS=3.12e-06 M=1 sca=1.01825
+ scb=8.55974e-05 scc=2.37716e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06
+ sa=1.2e-07 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M2@2 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.728e-13 PD=1.58e-06 PS=3.12e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06 sa=1.2e-07 sb=1.44e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/M2@3 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.728e-13 PD=1.58e-06 PS=3.12e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06 sa=1.2e-07 sb=1.44e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/M2@4 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.008e-13 PD=1.58e-06 PS=1.58e-06 M=1 sca=14.7929
+ scb=0.0126174 scc=0.00176209 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06
+ sa=5.6e-07 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M2@5 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.008e-13 PD=1.58e-06 PS=1.58e-06 M=1 sca=1.01825
+ scb=8.55974e-05 scc=2.37716e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06
+ sa=5.6e-07 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M2@6 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.008e-13 PD=1.58e-06 PS=1.58e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06 sa=5.6e-07 sb=1e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M2@7 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.008e-13 PD=1.58e-06 PS=1.58e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06 sa=5.6e-07 sb=1e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M2@8 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.008e-13 PD=1.58e-06 PS=1.58e-06 M=1 sca=14.7929
+ scb=0.0126174 scc=0.00176209 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06
+ sa=1e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M1@2 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.008e-13 PD=1.58e-06 PS=1.58e-06 M=1 sca=1.01825
+ scb=8.55974e-05 scc=2.37716e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06
+ sa=1e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M1@3 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.008e-13 PD=1.58e-06 PS=1.58e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06 sa=1e-06 sb=5.6e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M1@4 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.008e-13 PD=1.58e-06 PS=1.58e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06 sa=1e-06 sb=5.6e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M1@5 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.728e-13 PD=1.58e-06 PS=3.12e-06 M=1 sca=14.7929
+ scb=0.0126174 scc=0.00176209 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06
+ sa=1.44e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M1@6 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.728e-13 PD=1.58e-06 PS=3.12e-06 M=1 sca=1.01825
+ scb=8.55974e-05 scc=2.37716e-08 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06
+ sa=1.44e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/M1@7 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.728e-13 PD=1.58e-06 PS=3.12e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06 sa=1.44e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/M1@8 XI2/VBG XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=1.44e-06
+ AD=1.008e-13 AS=1.728e-13 PD=1.58e-06 PS=3.12e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.296e-06 sa=1.44e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XG2/M1 XI2/XI0/N3 XI2/VBP VDDHA_RX VDDHA_RX egpfet L=3e-07 W=8e-06
+ AD=5.6e-13 AS=9.6e-13 PD=8.14e-06 PS=1.624e-05 M=1 sca=4.68374 scb=0.00263327
+ scc=0.000317352 lpccnr=2.85e-07 covpccnr=0 wrxcnr=7.2e-06 sa=1.2e-07
+ sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/XG2/M2 XI2/XI0/N3 XI2/XI0/PDB VDDHA_RX VDDHA_RX egpfet L=3e-07 W=8e-06
+ AD=5.6e-13 AS=9.6e-13 PD=8.14e-06 PS=1.624e-05 M=1 sca=5.79873 scb=0.00379596
+ scc=0.000321345 lpccnr=2.85e-07 covpccnr=0 wrxcnr=7.2e-06 sa=5.6e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/XG2/M4 XI2/XI0/XG2/N1 XI2/XI0/PDB VSSA_RX VSSA_RX egnfet L=8e-06
+ W=4.2e-07 AD=5.04e-14 AS=5.04e-14 PD=1.08e-06 PS=1.08e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=7.215e-06 covpccnr=0 wrxcnr=3.78e-07 sa=1.2e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XG2/M3 XI2/XI0/N3 XI2/VBP XI2/XI0/XG2/N1 VSSA_RX egnfet L=8e-06
+ W=4.2e-07 AD=5.04e-14 AS=5.04e-14 PD=1.08e-06 PS=1.08e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=7.215e-06 covpccnr=0 wrxcnr=3.78e-07 sa=1.2e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/RRD4@2 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 20258.9 M=1 w=1e-06
+ l=3.326e-05   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/RRD4 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 20258.9 M=1 w=1e-06
+ l=3.326e-05   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/RRD3@2 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 5600 M=1 w=1e-06 l=9.1e-06  
+ bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/RRD3 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 5600 M=1 w=1e-06 l=9.1e-06  
+ bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR2/RR1 X290/X12/X50/X4/noxref_5 XI2/VBG VDDHA_RX opppcres 2784.36 M=1
+ w=2e-06 l=9.1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR2/RR2 X290/X12/X50/X4/noxref_5 X290/X12/X50/X4/noxref_6 VDDHA_RX
+ opppcres 2784.36 M=1 w=2e-06 l=9.1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR2/RR3 X290/X12/X50/X4/noxref_7 X290/X12/X50/X4/noxref_6 VDDHA_RX
+ opppcres 2784.36 M=1 w=2e-06 l=9.1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR2/RR4 X290/X12/X50/X4/noxref_7 X290/X12/X50/X4/noxref_8 VDDHA_RX
+ opppcres 2784.36 M=1 w=2e-06 l=9.1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR2/RR5 XI2/XI0/INP X290/X12/X50/X4/noxref_8 VDDHA_RX opppcres 2784.36
+ M=1 w=2e-06 l=9.1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR1/RR1 X290/X12/X50/X5/noxref_5 XI2/VBG VDDHA_RX opppcres 2784.36 M=1
+ w=2e-06 l=9.1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR1/RR2 X290/X12/X50/X5/noxref_5 X290/X12/X50/X5/noxref_6 VDDHA_RX
+ opppcres 2784.36 M=1 w=2e-06 l=9.1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR1/RR3 X290/X12/X50/X5/noxref_7 X290/X12/X50/X5/noxref_6 VDDHA_RX
+ opppcres 2784.36 M=1 w=2e-06 l=9.1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR1/RR4 X290/X12/X50/X5/noxref_7 X290/X12/X50/X5/noxref_8 VDDHA_RX
+ opppcres 2784.36 M=1 w=2e-06 l=9.1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR1/RR5 XI2/XI0/INN X290/X12/X50/X5/noxref_8 VDDHA_RX opppcres 2784.36
+ M=1 w=2e-06 l=9.1e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIRC/RR1 X290/X12/X50/noxref_8 XI2/VBG VDDHA_RX opppcres 968.268 M=1
+ w=2e-06 l=3.08e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIRC/RR2 X290/X12/X50/noxref_8 XI2/XI0/N2 VDDHA_RX opppcres 968.268 M=1
+ w=2e-06 l=3.08e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR3/RR1 X290/X12/X50/noxref_9 XI2/XI0/INP VDDHA_RX opppcres 1043.69
+ M=1 w=2e-06 l=3.33e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XIR3/RR2 X290/X12/X50/noxref_9 XI2/XI0/N1 VDDHA_RX opppcres 1043.69 M=1
+ w=2e-06 l=3.33e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/XOP/M18 XI2/XI0/XOP/N8 XI2/XI0/XOP/N8 XI2/XI0/XOP/N1N22 VSSA_RX egnfet
+ L=6e-07 W=6.2e-07 AD=4.34e-14 AS=7.44e-14 PD=7.6e-07 PS=1.48e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=1.2e-07 sb=8.6e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M16 XI2/XI0/XOP/N1N22 XI2/XI0/XOP/N8 VSSA_RX VSSA_RX egnfet
+ L=1.2e-06 W=5e-07 AD=6e-14 AS=6e-14 PD=1.24e-06 PS=1.24e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.095e-06 covpccnr=0 wrxcnr=4.5e-07 sa=1.2e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M18@2 XI2/XI0/XOP/N8 XI2/XI0/XOP/N8 XI2/XI0/XOP/N1N22 VSSA_RX
+ egnfet L=6e-07 W=6.2e-07 AD=4.34e-14 AS=7.44e-14 PD=7.6e-07 PS=1.48e-06 M=1
+ sca=0 scb=0 scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07 sa=8.6e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M15 XI2/XI0/XOP/N1N24 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=7.44e-14 PD=7.6e-07 PS=1.48e-06 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=1.2e-07 sb=8.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M17 XI2/XI0/XOP/N7 XI2/XI0/XOP/N8 XI2/XI0/XOP/N1N24 VSSA_RX egnfet
+ L=6e-07 W=1.54e-06 AD=1.078e-13 AS=1.848e-13 PD=1.68e-06 PS=3.32e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06 sa=1.2e-07 sb=8.6e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M15@2 XI2/XI0/XOP/N1N24 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet
+ L=6e-07 W=6.2e-07 AD=4.34e-14 AS=7.44e-14 PD=7.6e-07 PS=1.48e-06 M=1
+ sca=0.975587 scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0
+ wrxcnr=5.58e-07 sa=8.6e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M17@2 XI2/XI0/XOP/N7 XI2/XI0/XOP/N8 XI2/XI0/XOP/N1N24 VSSA_RX
+ egnfet L=6e-07 W=1.54e-06 AD=1.078e-13 AS=1.848e-13 PD=1.68e-06 PS=3.32e-06
+ M=1 sca=0 scb=0 scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06 sa=8.6e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M11 XI2/XI0/XOP/N1 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=7.44e-14 PD=7.6e-07 PS=1.48e-06 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M11@6 XI2/XI0/XOP/N1 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=4.34e-14 PD=7.6e-07 PS=7.6e-07 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=8.6e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M11@5 XI2/XI0/XOP/N1 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=4.34e-14 PD=7.6e-07 PS=7.6e-07 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=1.6e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M11@4 XI2/XI0/XOP/N1 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=4.34e-14 PD=7.6e-07 PS=7.6e-07 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=2.0083e-06 sb=1.6e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M11@3 XI2/XI0/XOP/N1 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=4.34e-14 PD=7.6e-07 PS=7.6e-07 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=2.0083e-06 sb=8.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M11@2 XI2/XI0/XOP/N1 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=7.44e-14 PD=7.6e-07 PS=1.48e-06 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M13 XI2/XI0/XOP/N7 XI2/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M12 XI2/XI0/XOP/N2 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=7.44e-14 PD=7.6e-07 PS=1.48e-06 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M12@6 XI2/XI0/XOP/N2 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=4.34e-14 PD=7.6e-07 PS=7.6e-07 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=8.6e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M12@5 XI2/XI0/XOP/N2 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=4.34e-14 PD=7.6e-07 PS=7.6e-07 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=1.6e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M12@4 XI2/XI0/XOP/N2 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=4.34e-14 PD=7.6e-07 PS=7.6e-07 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=2.0083e-06 sb=1.6e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M12@3 XI2/XI0/XOP/N2 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=4.34e-14 PD=7.6e-07 PS=7.6e-07 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=2.0083e-06 sb=8.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M12@2 XI2/XI0/XOP/N2 XI2/XI0/XOP/N7 VSSA_RX VSSA_RX egnfet L=6e-07
+ W=6.2e-07 AD=4.34e-14 AS=7.44e-14 PD=7.6e-07 PS=1.48e-06 M=1 sca=0.975587
+ scb=4.61901e-05 scc=3.11883e-09 lpccnr=5.55e-07 covpccnr=0 wrxcnr=5.58e-07
+ sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M22 XI2/XI0/XOP/N1N21 XI2/XI0/XOP/N9 VDDHA_RX VDDHA_RX egpfet
+ L=4e-07 W=7.2e-07 AD=8.64e-14 AS=8.64e-14 PD=1.68e-06 PS=1.68e-06 M=1
+ sca=25.7732 scb=0.022048 scc=0.00349193 lpccnr=3.75e-07 covpccnr=0
+ wrxcnr=6.48e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M24 XI2/XI0/XOP/N9 XI2/XI0/XOP/N9 XI2/XI0/XOP/N1N21 VDDHA_RX egpfet
+ L=3e-07 W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1
+ sca=11.7371 scb=0.00975878 scc=0.00134975 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=1.692e-06 sa=1.2e-07 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M24@2 XI2/XI0/XOP/N9 XI2/XI0/XOP/N9 XI2/XI0/XOP/N1N21 VDDHA_RX
+ egpfet L=3e-07 W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1
+ sca=11.7371 scb=0.00975878 scc=0.00134975 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=1.692e-06 sa=5.6e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M23 XI2/XI0/XOP/N10 XI2/XI0/XOP/N9 XI2/XI0/XOP/N1N4 VDDHA_RX egpfet
+ L=3e-07 W=3.76e-06 AD=2.632e-13 AS=4.512e-13 PD=3.9e-06 PS=7.76e-06 M=1
+ sca=6.23441 scb=0.004892 scc=0.000674877 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.384e-06 sa=1.2e-07 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M21 XI2/XI0/XOP/N1N4 XI2/XI0/XOP/N10 VDDHA_RX VDDHA_RX egpfet
+ L=3e-07 W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.2e-07 sb=5.6e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M23@2 XI2/XI0/XOP/N10 XI2/XI0/XOP/N9 XI2/XI0/XOP/N1N4 VDDHA_RX
+ egpfet L=3e-07 W=3.76e-06 AD=2.632e-13 AS=4.512e-13 PD=3.9e-06 PS=7.76e-06 M=1
+ sca=6.23441 scb=0.004892 scc=0.000674877 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.384e-06 sa=5.6e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M21@2 XI2/XI0/XOP/N1N4 XI2/XI0/XOP/N10 VDDHA_RX VDDHA_RX egpfet
+ L=3e-07 W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=5.6e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M19 XI2/XI0/XOP/N8 XI2/XI0/XOP/N10 VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.2e-07 sb=5.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M19@2 XI2/XI0/XOP/N8 XI2/XI0/XOP/N10 VDDHA_RX VDDHA_RX egpfet
+ L=3e-07 W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=5.6e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M20 XI2/XI0/XOP/N7 XI2/XI0/XOP/N10 VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.2e-07 sb=5.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M20@2 XI2/XI0/XOP/N7 XI2/XI0/XOP/N10 VDDHA_RX VDDHA_RX egpfet
+ L=3e-07 W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=5.6e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M7 XI2/XI0/XOP/N6 XI2/XI0/XOP/N9 XI2/XI0/XOP/N4 VDDHA_RX egpfet
+ L=3e-07 W=3.76e-06 AD=2.632e-13 AS=4.512e-13 PD=3.9e-06 PS=7.76e-06 M=1
+ sca=6.23441 scb=0.004892 scc=0.000674877 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.384e-06 sa=1.2e-07 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M7@4 XI2/XI0/XOP/N6 XI2/XI0/XOP/N9 XI2/XI0/XOP/N4 VDDHA_RX egpfet
+ L=3e-07 W=3.76e-06 AD=2.632e-13 AS=2.632e-13 PD=3.9e-06 PS=3.9e-06 M=1
+ sca=6.23441 scb=0.004892 scc=0.000674877 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.384e-06 sa=5.6e-07 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M7@3 XI2/XI0/XOP/N6 XI2/XI0/XOP/N9 XI2/XI0/XOP/N4 VDDHA_RX egpfet
+ L=3e-07 W=3.76e-06 AD=2.632e-13 AS=2.632e-13 PD=3.9e-06 PS=3.9e-06 M=1
+ sca=6.23441 scb=0.004892 scc=0.000674877 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.384e-06 sa=1e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M7@2 XI2/XI0/XOP/N6 XI2/XI0/XOP/N9 XI2/XI0/XOP/N4 VDDHA_RX egpfet
+ L=3e-07 W=3.76e-06 AD=2.632e-13 AS=4.512e-13 PD=3.9e-06 PS=7.76e-06 M=1
+ sca=6.23441 scb=0.004892 scc=0.000674877 lpccnr=2.85e-07 covpccnr=0
+ wrxcnr=3.384e-06 sa=1.44e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/MD VDDHA_RX VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=4e-06
+ AD=4.8e-13 AS=4.8e-13 PD=8.24e-06 PS=8.24e-06 M=1 sca=5.88235 scb=0.00459849
+ scc=0.000634384 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M1 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=4.8e-13 PD=4.14e-06 PS=8.24e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M1@16 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=5.4e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M1@15 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=9.6e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M1@14 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.38e-06 sb=1.8e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M1@13 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.8e-06 sb=1.38e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M1@12 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=9.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M1@11 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M1@10 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=4.8e-13 PD=4.14e-06 PS=8.24e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M2 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=4.8e-13 PD=4.14e-06 PS=8.24e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M2@16 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=5.4e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M2@15 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=9.6e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M2@14 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.38e-06 sb=1.8e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M2@13 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=1.8e-06 sb=1.38e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M2@12 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=9.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M2@11 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=5.4e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M2@10 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=4.8e-13 PD=4.14e-06 PS=8.24e-06 M=1
+ sca=5.88235 scb=0.00459849 scc=0.000634384 lpccnr=2.67e-07 covpccnr=0
+ wrxcnr=3.6e-06 sa=2.0083e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/MD@4 VDDHA_RX VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=4e-06
+ AD=4.8e-13 AS=4.8e-13 PD=8.24e-06 PS=8.24e-06 M=1 sca=5.88235 scb=0.00459849
+ scc=0.000634384 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M8 XI2/VBP XI2/XI0/XOP/N9 XI2/XI0/XOP/N5 VDDHA_RX egpfet L=3e-07
+ W=3.76e-06 AD=2.632e-13 AS=4.512e-13 PD=3.9e-06 PS=7.76e-06 M=1 sca=6.23441
+ scb=0.004892 scc=0.000674877 lpccnr=2.85e-07 covpccnr=0 wrxcnr=3.384e-06
+ sa=1.2e-07 sb=1.44e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M8@4 XI2/VBP XI2/XI0/XOP/N9 XI2/XI0/XOP/N5 VDDHA_RX egpfet L=3e-07
+ W=3.76e-06 AD=2.632e-13 AS=2.632e-13 PD=3.9e-06 PS=3.9e-06 M=1 sca=6.23441
+ scb=0.004892 scc=0.000674877 lpccnr=2.85e-07 covpccnr=0 wrxcnr=3.384e-06
+ sa=5.6e-07 sb=1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M8@3 XI2/VBP XI2/XI0/XOP/N9 XI2/XI0/XOP/N5 VDDHA_RX egpfet L=3e-07
+ W=3.76e-06 AD=2.632e-13 AS=2.632e-13 PD=3.9e-06 PS=3.9e-06 M=1 sca=6.23441
+ scb=0.004892 scc=0.000674877 lpccnr=2.85e-07 covpccnr=0 wrxcnr=3.384e-06
+ sa=1e-06 sb=5.6e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M8@2 XI2/VBP XI2/XI0/XOP/N9 XI2/XI0/XOP/N5 VDDHA_RX egpfet L=3e-07
+ W=3.76e-06 AD=2.632e-13 AS=4.512e-13 PD=3.9e-06 PS=7.76e-06 M=1 sca=6.23441
+ scb=0.004892 scc=0.000674877 lpccnr=2.85e-07 covpccnr=0 wrxcnr=3.384e-06
+ sa=1.44e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M9 XI2/XI0/XOP/N6 XI2/XI0/XOP/N8 XI2/XI0/XOP/N1 VSSA_RX egnfet
+ L=6e-07 W=1.54e-06 AD=1.078e-13 AS=1.848e-13 PD=1.68e-06 PS=3.32e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M9@4 XI2/XI0/XOP/N6 XI2/XI0/XOP/N8 XI2/XI0/XOP/N1 VSSA_RX egnfet
+ L=6e-07 W=1.54e-06 AD=1.078e-13 AS=1.078e-13 PD=1.68e-06 PS=1.68e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06 sa=8.6e-07 sb=1.6e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M9@3 XI2/XI0/XOP/N6 XI2/XI0/XOP/N8 XI2/XI0/XOP/N1 VSSA_RX egnfet
+ L=6e-07 W=1.54e-06 AD=1.078e-13 AS=1.078e-13 PD=1.68e-06 PS=1.68e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06 sa=1.6e-06 sb=8.6e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M9@2 XI2/XI0/XOP/N6 XI2/XI0/XOP/N8 XI2/XI0/XOP/N1 VSSA_RX egnfet
+ L=6e-07 W=1.54e-06 AD=1.078e-13 AS=1.848e-13 PD=1.68e-06 PS=3.32e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M5 XI2/XI0/XOP/N4 XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.2e-07 sb=1.44e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M5@4 XI2/XI0/XOP/N4 XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.88e-06 AD=1.316e-13 AS=1.316e-13 PD=2.02e-06 PS=2.02e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=5.6e-07 sb=1e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M5@3 XI2/XI0/XOP/N4 XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.88e-06 AD=1.316e-13 AS=1.316e-13 PD=2.02e-06 PS=2.02e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1e-06 sb=5.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M5@2 XI2/XI0/XOP/N4 XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.44e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/MD@3 VDDHA_RX VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=4e-06
+ AD=4.8e-13 AS=4.8e-13 PD=8.24e-06 PS=8.24e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M1@9 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=4.8e-13 PD=4.14e-06 PS=8.24e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.2e-07 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M1@8 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=5.4e-07 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M1@7 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=9.6e-07 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M1@6 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.38e-06 sb=1.8e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M1@5 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.8e-06 sb=1.38e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M1@4 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=9.6e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M3 XI2/XI0/XOP/N3 XI2/XI0/XOP/N10 VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.2e-07 sb=5.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M1@3 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=5.4e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M1@2 XI2/XI0/XOP/N1 XI2/XI0/INP XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=4.8e-13 PD=4.14e-06 PS=8.24e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M3@4 XI2/XI0/XOP/N3 XI2/XI0/XOP/N10 VDDHA_RX VDDHA_RX egpfet
+ L=3e-07 W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=5.6e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M10 XI2/VBP XI2/XI0/XOP/N8 XI2/XI0/XOP/N2 VSSA_RX egnfet L=6e-07
+ W=1.54e-06 AD=1.078e-13 AS=1.848e-13 PD=1.68e-06 PS=3.32e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06 sa=1.2e-07 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M10@4 XI2/VBP XI2/XI0/XOP/N8 XI2/XI0/XOP/N2 VSSA_RX egnfet L=6e-07
+ W=1.54e-06 AD=1.078e-13 AS=1.078e-13 PD=1.68e-06 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06 sa=8.6e-07 sb=1.6e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M10@3 XI2/VBP XI2/XI0/XOP/N8 XI2/XI0/XOP/N2 VSSA_RX egnfet L=6e-07
+ W=1.54e-06 AD=1.078e-13 AS=1.078e-13 PD=1.68e-06 PS=1.68e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06 sa=1.6e-06 sb=8.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M10@2 XI2/VBP XI2/XI0/XOP/N8 XI2/XI0/XOP/N2 VSSA_RX egnfet L=6e-07
+ W=1.54e-06 AD=1.078e-13 AS=1.848e-13 PD=1.68e-06 PS=3.32e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=5.55e-07 covpccnr=0 wrxcnr=1.386e-06 sa=2.0083e-06 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M6 XI2/XI0/XOP/N5 XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.2e-07 sb=1.44e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M6@4 XI2/XI0/XOP/N5 XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.88e-06 AD=1.316e-13 AS=1.316e-13 PD=2.02e-06 PS=2.02e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=5.6e-07 sb=1e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M6@3 XI2/XI0/XOP/N5 XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.88e-06 AD=1.316e-13 AS=1.316e-13 PD=2.02e-06 PS=2.02e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1e-06 sb=5.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M6@2 XI2/XI0/XOP/N5 XI2/XI0/XOP/N6 VDDHA_RX VDDHA_RX egpfet L=3e-07
+ W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.44e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/MD@2 VDDHA_RX VDDHA_RX VDDHA_RX VDDHA_RX egpfet L=2.8e-07 W=4e-06
+ AD=4.8e-13 AS=4.8e-13 PD=8.24e-06 PS=8.24e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M2@9 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=4.8e-13 PD=4.14e-06 PS=8.24e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.2e-07 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M2@8 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=5.4e-07 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M2@7 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=9.6e-07 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M2@6 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.38e-06 sb=1.8e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M2@5 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=1.8e-06 sb=1.38e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M2@4 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=9.6e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M3@3 XI2/XI0/XOP/N3 XI2/XI0/XOP/N10 VDDHA_RX VDDHA_RX egpfet
+ L=3e-07 W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=1.2e-07 sb=5.6e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M2@3 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=2.8e-13 PD=4.14e-06 PS=4.14e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=5.4e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M2@2 XI2/XI0/XOP/N2 XI2/XI0/INN XI2/XI0/XOP/N3 VDDHA_RX egpfet
+ L=2.8e-07 W=4e-06 AD=2.8e-13 AS=4.8e-13 PD=4.14e-06 PS=8.24e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.67e-07 covpccnr=0 wrxcnr=3.6e-06 sa=2.0083e-06 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M3@2 XI2/XI0/XOP/N3 XI2/XI0/XOP/N10 VDDHA_RX VDDHA_RX egpfet
+ L=3e-07 W=1.88e-06 AD=1.316e-13 AS=2.256e-13 PD=2.02e-06 PS=4e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=2.85e-07 covpccnr=0 wrxcnr=1.692e-06 sa=5.6e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/M26 XI2/XI0/XOP/N9 XI2/XI0/XOP/N14 VSSA_RX VSSA_RX egnfet L=7e-07
+ W=4.6e-07 AD=3.22e-14 AS=5.52e-14 PD=6e-07 PS=1.16e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=1.2e-07 sb=9.6e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M26@2 XI2/XI0/XOP/N9 XI2/XI0/XOP/N14 VSSA_RX VSSA_RX egnfet L=7e-07
+ W=4.6e-07 AD=3.22e-14 AS=5.52e-14 PD=6e-07 PS=1.16e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=9.6e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M25 XI2/XI0/XOP/N10 XI2/XI0/XOP/N14 VSSA_RX VSSA_RX egnfet L=7e-07
+ W=4.6e-07 AD=3.22e-14 AS=5.52e-14 PD=6e-07 PS=1.16e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=1.2e-07 sb=9.6e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/M25@2 XI2/XI0/XOP/N10 XI2/XI0/XOP/N14 VSSA_RX VSSA_RX egnfet
+ L=7e-07 W=4.6e-07 AD=3.22e-14 AS=5.52e-14 PD=6e-07 PS=1.16e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=9.6e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/CC0 XI2/VBP XI2/XI0/N2 VSSA_RX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI0/CC1 XI2/XI0/N2 XI2/VBP VSSA_RX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI0/CC2 XI2/VBP XI2/XI0/N2 VSSA_RX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI0/CC3 XI2/XI0/N2 XI2/VBP VSSA_RX vncap  botcap=0 botlev=17 setind=-2
+ toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI0/Q21 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q22 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q23 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q24 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q25 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q26 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q27 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q28 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q29 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q210 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q211 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q212 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q1 VSSA_RX VSSA_RX XI2/XI0/INN  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q213 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q214 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XXI2/XI0/Q215 VSSA_RX VSSA_RX XI2/XI0/N1  vpnp W=1e-05 L=1e-05 nf=1 nrep=1
+ sizedup=0
XX290/X12/X58/D0_noxref VSS XI2/XI0/XOP/XI0/N3 diodenwx  AREA=1.31355e-11
+ perim=1.451e-05 sizedup=0
XXI2/XI0/XOP/XI0/M6 XI2/XI0/XOP/N14 XI2/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M7 XI2/XI0/XOP/XI0/N4 XI2/PDI VSSA_RX VSSA_RX egnfet L=4.2e-07
+ W=2.5e-06 AD=3e-13 AS=3e-13 PD=5.24e-06 PS=5.24e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.93e-07 covpccnr=0 wrxcnr=2.25e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M8 XI2/XI0/XOP/XI0/N4 XI2/XI0/XOP/N14 VSSA_RX VSSA_RX egnfet
+ L=4.2e-07 W=2.5e-06 AD=3e-13 AS=3e-13 PD=5.24e-06 PS=5.24e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=3.93e-07 covpccnr=0 wrxcnr=2.25e-06 sa=1.2e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/XI0/M5 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/XI0/N4 VSSA_RX VSSA_RX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0
+ scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/XI0/X1I44/M0 XI2/XI0/XOP/XI0/TIEL XI2/XI0/XOP/XI0/X1I44/N1N50
+ VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06
+ PS=1.04e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M10 XI2/XI0/XOP/XI0/N4 XI2/XI0/XOP/N14 XI2/XI0/XOP/XI0/N1N5
+ VDDHA_RX egpfet L=2.5e-06 W=4.2e-07 AD=5.04e-14 AS=5.04e-14 PD=1.08e-06
+ PS=1.08e-06 M=1 sca=41.3582 scb=0.0318885 scc=0.00571618 lpccnr=2.265e-06
+ covpccnr=0 wrxcnr=3.78e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M10@2 XI2/XI0/XOP/XI0/N4 XI2/XI0/XOP/N14 XI2/XI0/XOP/XI0/N1N5
+ VDDHA_RX egpfet L=2.5e-06 W=4.2e-07 AD=5.04e-14 AS=5.04e-14 PD=1.08e-06
+ PS=1.08e-06 M=1 sca=9.94988 scb=0.00979913 scc=0.000251034 lpccnr=2.265e-06
+ covpccnr=0 wrxcnr=3.78e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M9 XI2/XI0/XOP/XI0/N1N5 XI2/PDI VDDHA_RX VDDHA_RX egpfet
+ L=2.5e-06 W=4.2e-07 AD=5.04e-14 AS=5.04e-14 PD=1.08e-06 PS=1.08e-06 M=1
+ sca=5.09368 scb=0.00317154 scc=0.00011934 lpccnr=2.265e-06 covpccnr=0
+ wrxcnr=3.78e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M9@2 XI2/XI0/XOP/XI0/N1N5 XI2/PDI VDDHA_RX VDDHA_RX egpfet
+ L=2.5e-06 W=4.2e-07 AD=5.04e-14 AS=5.04e-14 PD=1.08e-06 PS=1.08e-06 M=1
+ sca=4.04474 scb=0.00311197 scc=0.000119335 lpccnr=2.265e-06 covpccnr=0
+ wrxcnr=3.78e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M3 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/XI0/N2 VDDHA_RX VDDHA_RX
+ egpfet L=5.4e-07 W=1.2e-06 AD=8.4e-14 AS=1.44e-13 PD=1.34e-06 PS=2.64e-06 M=1
+ sca=5.29595 scb=0.00355861 scc=2.98846e-05 lpccnr=5.01e-07 covpccnr=0
+ wrxcnr=1.08e-06 sa=1.2e-07 sb=8e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M3@2 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/XI0/N2 VDDHA_RX VDDHA_RX
+ egpfet L=5.4e-07 W=1.2e-06 AD=8.4e-14 AS=1.44e-13 PD=1.34e-06 PS=2.64e-06 M=1
+ sca=22.2571 scb=0.0220844 scc=0.00275492 lpccnr=5.01e-07 covpccnr=0
+ wrxcnr=1.08e-06 sa=8e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M4 XI2/XI0/XOP/N14 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/XI0/N3
+ XI2/XI0/XOP/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=8.4e-14 AS=1.44e-13
+ PD=1.34e-06 PS=2.64e-06 M=1 sca=27.3358 scb=0.0265429 scc=0.00265366
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/XI0/M4@8 XI2/XI0/XOP/N14 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/XI0/N3
+ XI2/XI0/XOP/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=8.4e-14 AS=1.44e-13
+ PD=1.34e-06 PS=2.64e-06 M=1 sca=15.6494 scb=0.0172079 scc=0.000712039
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/XI0/M4@7 XI2/XI0/XOP/N14 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/XI0/N3
+ XI2/XI0/XOP/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=8.4e-14 AS=8.4e-14
+ PD=1.34e-06 PS=1.34e-06 M=1 sca=22.1568 scb=0.0165232 scc=0.00211861
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=8e-07 sb=1.48e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M4@6 XI2/XI0/XOP/N14 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/XI0/N3
+ XI2/XI0/XOP/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=8.4e-14 AS=8.4e-14
+ PD=1.34e-06 PS=1.34e-06 M=1 sca=10.4704 scb=0.00718825 scc=0.00017699
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=8e-07 sb=1.48e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M4@5 XI2/XI0/XOP/N14 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/XI0/N3
+ XI2/XI0/XOP/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=8.4e-14 AS=8.4e-14
+ PD=1.34e-06 PS=1.34e-06 M=1 sca=22.1568 scb=0.0165232 scc=0.00211861
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.48e-06 sb=8e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M4@4 XI2/XI0/XOP/N14 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/XI0/N3
+ XI2/XI0/XOP/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=8.4e-14 AS=8.4e-14
+ PD=1.34e-06 PS=1.34e-06 M=1 sca=10.4704 scb=0.00718825 scc=0.00017699
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=1.48e-06 sb=8e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/M4@3 XI2/XI0/XOP/N14 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/XI0/N3
+ XI2/XI0/XOP/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=8.4e-14 AS=1.44e-13
+ PD=1.34e-06 PS=2.64e-06 M=1 sca=27.3358 scb=0.0265429 scc=0.00265366
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/XI0/M4@2 XI2/XI0/XOP/N14 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/XI0/N3
+ XI2/XI0/XOP/XI0/N3 egpfet L=5.4e-07 W=1.2e-06 AD=8.4e-14 AS=1.44e-13
+ PD=1.34e-06 PS=2.64e-06 M=1 sca=15.6494 scb=0.0172079 scc=0.000712039
+ lpccnr=5.01e-07 covpccnr=0 wrxcnr=1.08e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/XI0/MR XI2/XI0/XOP/XI0/N3 XI2/XI0/XOP/XI0/TIEL VDDHA_RX VDDHA_RX
+ egpfet L=8e-07 W=5.2e-07 AD=6.24e-14 AS=6.24e-14 PD=1.28e-06 PS=1.28e-06 M=1
+ sca=48.5924 scb=0.0434689 scc=0.00660393 lpccnr=7.35e-07 covpccnr=0
+ wrxcnr=4.68e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI0/XOP/XI0/X1I44/M1 XI2/XI0/XOP/XI0/X1I44/N1N50
+ XI2/XI0/XOP/XI0/X1I44/N1N50 VDDHA_RX VDDHA_RX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=40.863 scb=0.0302947
+ scc=0.00581109 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/XI0/M1 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/N14 VSSA_RX VSSA_RX egnfet
+ L=7e-07 W=4.6e-07 AD=3.22e-14 AS=5.52e-14 PD=6e-07 PS=1.16e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=1.2e-07 sb=9.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/XI0/M1@2 XI2/XI0/XOP/XI0/N2 XI2/XI0/XOP/N14 VSSA_RX VSSA_RX egnfet
+ L=7e-07 W=4.6e-07 AD=3.22e-14 AS=5.52e-14 PD=6e-07 PS=1.16e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=9.6e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/XI0/M2 XI2/XI0/XOP/N14 XI2/XI0/XOP/N14 VSSA_RX VSSA_RX egnfet
+ L=7e-07 W=4.6e-07 AD=3.22e-14 AS=5.52e-14 PD=6e-07 PS=1.16e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=1.2e-07 sb=9.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI0/XOP/XI0/M2@2 XI2/XI0/XOP/N14 XI2/XI0/XOP/N14 VSSA_RX VSSA_RX egnfet
+ L=7e-07 W=4.6e-07 AD=3.22e-14 AS=5.52e-14 PD=6e-07 PS=1.16e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=6.45e-07 covpccnr=0 wrxcnr=4.14e-07 sa=9.6e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XX290/X13/D0_noxref VSS VDDHA_RX diodenwx  AREA=4.35278e-10 perim=0.00010032
+ sizedup=0
XX290/X13/D1_noxref VSS VDDHA_RX diodenwx  AREA=4.31842e-10 perim=0.00010575
+ sizedup=0
XXI2/XI1/X2I178/M1 XI2/XI1/TIEH5 XI2/XI1/X2I178/N1N42 VDDHA_RX VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=38.4615 scb=0.0292734 scc=0.00580942 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I176/M1 XI2/XI1/TIEH4 XI2/XI1/X2I176/N1N42 VDDHA_RX VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=39.7843 scb=0.02942 scc=0.00580945 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I174/M1 XI2/XI1/TIEH3 XI2/XI1/X2I174/N1N42 VDDHA_RX VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=41.548
+ scb=0.0311992 scc=0.00581613 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I171/M1 XI2/XI1/TIEH2 XI2/XI1/X2I171/N1N42 VDDHA_RX VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=52.3504 scb=0.0474888 scc=0.00707531 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XIRZ/RR1 XI2/XI1/VBP X290/X13/X6/noxref_30 VDDHA_RX opppcres 2090.5 M=1
+ w=2e-06 l=6.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/XIRZ/RR2 XI2/XI1/N1N209 X290/X13/X6/noxref_30 VDDHA_RX opppcres 2090.5
+ M=1 w=2e-06 l=6.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/M17 XI2/XI1/PDB XI2/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M8 XI2/N1N12 XI2/PDI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X1I241/M0 XI2/XI1/X1I241/N1N42 XI2/XI1/X1I241/N1N42 VSSA_RX VSSA_RX
+ egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M18E IBTX2 XI2/PDTXI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG9/M2 XI2/XI1/N2N116 XI2/CAI0 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06 PS=3.04e-06 M=1 sca=20.5863
+ scb=0.0188352 scc=0.00189527 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG9/M1 XI2/XI1/N2N116 XI2/XI1/PDTXB VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06 PS=3.04e-06 M=1 sca=18.5161
+ scb=0.0152985 scc=0.00182278 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M5 XI2/XI1/VBP XI2/XI1/N2 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=11.7416 scb=0.00859489
+ scc=0.00105884 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/XG10/M1 XI2/XI1/S0 XI2/XI1/N2N116 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=16.4041
+ scb=0.0130724 scc=0.00181242 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M5@4 XI2/XI1/VBP XI2/XI1/N2 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=10.8015
+ scb=0.00783256 scc=0.00105735 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=6.1e-07 sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M5@3 XI2/XI1/VBP XI2/XI1/N2 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=10.3381
+ scb=0.00769091 scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=1.1e-06 sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG11/M1 XI2/XI1/S0B XI2/XI1/S0 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=15.1515
+ scb=0.0129539 scc=0.00181241 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M5@2 XI2/XI1/VBP XI2/XI1/N2 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396
+ scb=0.00766114 scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=1.59e-06 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I71/M2 XI2/XI1/VBP XI2/XI1/S0B XI2/XI1/N2N77 VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=38.4615
+ scb=0.0292734 scc=0.00580942 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I71/M4 XI2/XI1/N2N77 XI2/XI1/S0 XI2/XI1/TIEH5 VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=38.4615
+ scb=0.0292734 scc=0.00580942 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10H IBTX2 XI2/XI1/N2N77 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10H@6 IBTX2 XI2/XI1/N2N77 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=6.1e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10H@5 IBTX2 XI2/XI1/N2N77 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10H@4 IBTX2 XI2/XI1/N2N77 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06
+ sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M4 XI2/XI1/N2 XI2/XI1/N2 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10H@3 IBTX2 XI2/XI1/N2N77 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M4@4 XI2/XI1/N2 XI2/XI1/N2 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=6.1e-07 sb=1.1e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10H@2 IBTX2 XI2/XI1/N2N77 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M4@3 XI2/XI1/N2 XI2/XI1/N2 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06 sb=6.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M4@2 XI2/XI1/N2 XI2/XI1/N2 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M16 XI2/XI1/PDB XI2/PDI VDDHA_RX VDDHA_RX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=31.2344 scb=0.0274471
+ scc=0.00468985 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M9 XI2/XI1/VBP XI2/XI1/PDB VDDHA_RX VDDHA_RX egpfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=2.57743 scb=0.00126348
+ scc=3.08066e-06 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M6 XI2/GMOUT XI2/XI1/VBP VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=8.01179 scb=0.00705084
+ scc=0.000849657 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M6@8 XI2/GMOUT XI2/XI1/VBP VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07 sb=1.59e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M6@7 XI2/GMOUT XI2/XI1/VBP VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=8.01179 scb=0.00705084
+ scc=0.000849657 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=6.1e-07
+ sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M6@6 XI2/GMOUT XI2/XI1/VBP VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=6.1e-07 sb=1.1e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M6@5 XI2/GMOUT XI2/XI1/VBP VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=8.01179 scb=0.00705084
+ scc=0.000849657 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06
+ sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M6@4 XI2/GMOUT XI2/XI1/VBP VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06 sb=6.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M6@3 XI2/GMOUT XI2/XI1/VBP VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=8.01179 scb=0.00705084
+ scc=0.000849657 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M6@2 XI2/GMOUT XI2/XI1/VBP VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I23/M2 XI2/XI1/VBP XI2/PDTXI XI2/XI1/N2N4 VDDHA_RX egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=38.4615
+ scb=0.0292734 scc=0.00580942 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I23/M4 XI2/XI1/N2N4 XI2/XI1/PDTXB XI2/XI1/TIEH2 VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=38.4615
+ scb=0.0292734 scc=0.00580942 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X1I241/M1 XI2/XI1/TIEH1 XI2/XI1/X1I241/N1N42 VDDHA_RX VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=114.438 scb=0.0900098 scc=0.017762 lpccnr=1.5e-07 covpccnr=0
+ wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1
+ p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10E IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=2.00435 scb=0.00117262
+ scc=1.24607e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10E@12 IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10E@11 IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=2.00435 scb=0.00117262
+ scc=1.24607e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=6.1e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10E@10 IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=6.1e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10E@9 IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=2.00435 scb=0.00117262
+ scc=1.24607e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10E@8 IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10E@7 IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=2.00435 scb=0.00117262
+ scc=1.24607e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06
+ sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10E@6 IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06
+ sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10E@5 IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=2.00435 scb=0.00117262
+ scc=1.24607e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10E@4 IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10E@3 IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=2.00435 scb=0.00117262
+ scc=1.24607e-05 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10E@2 IBTX2 XI2/XI1/N2N4 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/X2I23/M3 XI2/XI1/TIEH2 XI2/PDTXI XI2/XI1/N2N4 VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I23/M1 XI2/XI1/N2N4 XI2/XI1/PDTXB XI2/XI1/VBP VSSA_RX egnfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=4.1e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/XG1/M2 XI2/XI1/PDTXB XI2/PDTXI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M18D IBTX1 XI2/PDTXI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG1/M1 XI2/XI1/PDTXB XI2/PDTXI VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=15.1515
+ scb=0.0129539 scc=0.00181241 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I27/M2 XI2/XI1/VBP XI2/PDTXI XI2/XI1/N2N5 VDDHA_RX egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=38.4615
+ scb=0.0292734 scc=0.00580942 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I27/M4 XI2/XI1/N2N5 XI2/XI1/PDTXB XI2/XI1/TIEH2 VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=38.4615
+ scb=0.0292734 scc=0.00580942 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10D IBTX1 XI2/XI1/N2N5 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10D@10 IBTX1 XI2/XI1/N2N5 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=6.1e-07
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10D@9 IBTX1 XI2/XI1/N2N5 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10D@8 IBTX1 XI2/XI1/N2N5 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10D@7 IBTX1 XI2/XI1/N2N5 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10D@6 IBTX1 XI2/XI1/N2N5 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10D@5 IBTX1 XI2/XI1/N2N5 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=10.3437 scb=0.00774891
+ scc=0.00105732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10D@4 IBTX1 XI2/XI1/N2N5 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=11.191 scb=0.00815694
+ scc=0.00105784 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10D@3 IBTX1 XI2/XI1/N2N5 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=12.7412 scb=0.0101827
+ scc=0.00107638 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10D@2 IBTX1 XI2/XI1/N2N5 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=18.1291 scb=0.0184754
+ scc=0.00162359 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/X2I27/M3 XI2/XI1/TIEH2 XI2/PDTXI XI2/XI1/N2N5 VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I27/M1 XI2/XI1/N2N5 XI2/XI1/PDTXB XI2/XI1/VBP VSSA_RX egnfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=4.1e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/XG11/M2 XI2/XI1/S0B XI2/XI1/S0 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG10/M2 XI2/XI1/S0 XI2/XI1/N2N116 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG9/M3 XI2/XI1/N2N116 XI2/XI1/PDTXB XI2/XI1/XG9/N1 VSSA_RX egnfet
+ L=1.5e-07 W=8e-07 AD=9.6e-14 AS=5.6e-14 PD=1.84e-06 PS=9.4e-07 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=4.1e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/XG9/M4 XI2/XI1/XG9/N1 XI2/CAI0 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I71/M3 XI2/XI1/TIEH5 XI2/XI1/S0B XI2/XI1/N2N77 VSSA_RX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=4.1e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/X2I71/M1 XI2/XI1/N2N77 XI2/XI1/S0 XI2/XI1/VBP VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10F IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@25 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=6.59961
+ scb=0.00623493 scc=0.000619732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10F@24 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=6.1e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@23 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=6.59961
+ scb=0.00623493 scc=0.000619732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=6.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10F@22 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@21 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=6.59961
+ scb=0.00623493 scc=0.000619732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=1.1e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10F@20 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@19 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=6.59961
+ scb=0.00623493 scc=0.000619732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=1.59e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10F@18 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@17 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=6.59961
+ scb=0.00623493 scc=0.000619732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10F@16 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@15 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=6.59961
+ scb=0.00623493 scc=0.000619732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10F@14 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@13 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=6.59961
+ scb=0.00623493 scc=0.000619732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=2.0083e-06 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10F@12 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@11 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=6.59961
+ scb=0.00623493 scc=0.000619732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=2.0083e-06 sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10F@10 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=2.0083e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@9 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=6.59961 scb=0.00623493
+ scc=0.000619732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10F@8 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@7 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=6.59961 scb=0.00623493
+ scc=0.000619732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10F@6 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=1.59e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@5 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=2.88e-13 AS=1.68e-13 PD=5.04e-06 PS=2.54e-06 M=1 sca=6.59961 scb=0.00623493
+ scc=0.000619732 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10F@4 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=1.1e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@3 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=6.1e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10F@2 IBTX2 XI2/XI1/N2N42 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/X2I47/M4 XI2/XI1/N2N42 XI2/XI1/S2 XI2/XI1/TIEH3 VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=24.3167
+ scb=0.0247876 scc=0.00343783 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I47/M2 XI2/XI1/VBP XI2/XI1/S2B XI2/XI1/N2N42 VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=24.3167
+ scb=0.0247876 scc=0.00343783 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG5/M1 XI2/XI1/S2B XI2/XI1/S2 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=10.3816
+ scb=0.0105595 scc=0.00106234 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG4/M1 XI2/XI1/S2 XI2/XI1/N2N95 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=10.3816
+ scb=0.0105595 scc=0.00106234 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG3/M1 XI2/XI1/N2N95 XI2/XI1/PDTXB VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06 PS=3.04e-06 M=1 sca=10.3816
+ scb=0.0105595 scc=0.00106234 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG3/M2 XI2/XI1/N2N95 XI2/CAI2 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06 PS=3.04e-06 M=1 sca=10.3816
+ scb=0.0105595 scc=0.00106234 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG5/M2 XI2/XI1/S2B XI2/XI1/S2 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG4/M2 XI2/XI1/S2 XI2/XI1/N2N95 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG3/M3 XI2/XI1/N2N95 XI2/XI1/PDTXB XI2/XI1/XG3/N1 VSSA_RX egnfet
+ L=1.5e-07 W=8e-07 AD=9.6e-14 AS=5.6e-14 PD=1.84e-06 PS=9.4e-07 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=4.1e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/XG3/M4 XI2/XI1/XG3/N1 XI2/CAI2 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I47/M3 XI2/XI1/TIEH3 XI2/XI1/S2B XI2/XI1/N2N42 VSSA_RX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=4.1e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/X2I47/M1 XI2/XI1/N2N42 XI2/XI1/S2 XI2/XI1/VBP VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG0/M2 XI2/XI1/PDRXB XI2/PDRXI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M18 IBRX1 XI2/PDRXI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07 AD=4.8e-14
+ AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0 lpccnr=1.5e-07
+ covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M18B IBRX2 XI2/PDRXI VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG0/M1 XI2/XI1/PDRXB XI2/PDRXI VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=15.1515
+ scb=0.0129539 scc=0.00181241 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X1I82/M2 XI2/XI1/VBP XI2/PDRXI XI2/XI1/N1N83 VDDHA_RX egpfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=38.4615
+ scb=0.0292734 scc=0.00580942 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X1I82/M4 XI2/XI1/N1N83 XI2/XI1/PDRXB XI2/XI1/TIEH1 VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=38.4615
+ scb=0.0292734 scc=0.00580942 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10 IBRX1 XI2/XI1/N1N83 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10@4 IBRX1 XI2/XI1/N1N83 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=6.1e-07 sb=1.1e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10@3 IBRX1 XI2/XI1/N1N83 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06 sb=6.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10@2 IBRX1 XI2/XI1/N1N83 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10B IBRX2 XI2/XI1/N1N83 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10B@4 IBRX2 XI2/XI1/N1N83 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=6.1e-07 sb=1.1e-06
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10B@3 IBRX2 XI2/XI1/N1N83 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06 sb=6.1e-07
+ sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10B@2 IBRX2 XI2/XI1/N1N83 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/X1I82/M3 XI2/XI1/TIEH1 XI2/PDRXI XI2/XI1/N1N83 VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X1I82/M1 XI2/XI1/N1N83 XI2/XI1/PDRXB XI2/XI1/VBP VSSA_RX egnfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=4.1e-07 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/XG6/M2 XI2/XI1/N2N102 XI2/CAI1 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06 PS=3.04e-06 M=1 sca=15.1515
+ scb=0.0129539 scc=0.00181241 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG6/M1 XI2/XI1/N2N102 XI2/XI1/PDTXB VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=9.8e-14 AS=1.68e-13 PD=1.54e-06 PS=3.04e-06 M=1 sca=15.1515
+ scb=0.0129539 scc=0.00181241 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG7/M1 XI2/XI1/S1 XI2/XI1/N2N102 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=15.1515
+ scb=0.0129539 scc=0.00181241 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG8/M1 XI2/XI1/S1B XI2/XI1/S1 VDDHA_RX VDDHA_RX egpfet L=1.5e-07
+ W=1.4e-06 AD=1.68e-13 AS=1.68e-13 PD=3.04e-06 PS=3.04e-06 M=1 sca=15.1515
+ scb=0.0129539 scc=0.00181241 lpccnr=1.5e-07 covpccnr=0 wrxcnr=1.26e-06
+ sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I60/M2 XI2/XI1/VBP XI2/XI1/S1B XI2/XI1/N2N69 VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=38.4615
+ scb=0.0292734 scc=0.00580942 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=1.2e-07 sb=4.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I60/M4 XI2/XI1/N2N69 XI2/XI1/S1 XI2/XI1/TIEH4 VDDHA_RX egpfet
+ L=1.5e-07 W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=38.4615
+ scb=0.0292734 scc=0.00580942 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07
+ sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10G IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10G@12 IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396
+ scb=0.00766114 scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=1.2e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10G@11 IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0
+ scc=0 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=6.1e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10G@10 IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07
+ W=2.4e-06 AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396
+ scb=0.00766114 scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06
+ sa=6.1e-07 sb=2.0083e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1
+ pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10G@9 IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06 sb=1.59e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10G@8 IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.1e-06
+ sb=1.59e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10G@7 IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06 sb=1.1e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M10G@6 IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=1.59e-06
+ sb=1.1e-06 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10G@5 IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=6.1e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10G@4 IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=1.68e-13 PD=2.54e-06 PS=2.54e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=6.1e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/M10G@3 IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M10G@2 IBTX2 XI2/XI1/N2N69 VDDHA_RX VDDHA_RX egpfet L=3.5e-07 W=2.4e-06
+ AD=1.68e-13 AS=2.88e-13 PD=2.54e-06 PS=5.04e-06 M=1 sca=9.43396 scb=0.00766114
+ scc=0.00105731 lpccnr=3.3e-07 covpccnr=0 wrxcnr=2.16e-06 sa=2.0083e-06
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/XG8/M2 XI2/XI1/S1B XI2/XI1/S1 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=4e-07
+ AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG7/M2 XI2/XI1/S1 XI2/XI1/N2N102 VSSA_RX VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XG6/M3 XI2/XI1/N2N102 XI2/XI1/PDTXB XI2/XI1/XG6/N1 VSSA_RX egnfet
+ L=1.5e-07 W=8e-07 AD=9.6e-14 AS=5.6e-14 PD=1.84e-06 PS=9.4e-07 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=1.2e-07 sb=4.1e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/XG6/M4 XI2/XI1/XG6/N1 XI2/CAI1 VSSA_RX VSSA_RX egnfet L=1.5e-07 W=8e-07
+ AD=5.6e-14 AS=9.6e-14 PD=9.4e-07 PS=1.84e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=7.2e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/X2I60/M3 XI2/XI1/TIEH4 XI2/XI1/S1B XI2/XI1/N2N69 VSSA_RX egnfet
+ L=1.5e-07 W=4e-07 AD=4.8e-14 AS=2.8e-14 PD=1.04e-06 PS=5.4e-07 M=1 sca=0 scb=0
+ scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07 sb=4.1e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/X2I60/M1 XI2/XI1/N2N69 XI2/XI1/S1 XI2/XI1/VBP VSSA_RX egnfet L=1.5e-07
+ W=4e-07 AD=2.8e-14 AS=4.8e-14 PD=5.4e-07 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=4.1e-07 sb=1.2e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M2 XI2/XI1/VBP XI2/VBG XI2/XI1/N1 VSSA_RX egnfet L=5e-07 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.65e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M3 XI2/XI1/N1 XI2/N1N12 VSSA_RX VSSA_RX egnfet L=7e-07 W=9e-07
+ AD=6.3e-14 AS=1.08e-13 PD=1.04e-06 PS=2.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=8.1e-07 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M2@4 XI2/XI1/VBP XI2/VBG XI2/XI1/N1 VSSA_RX egnfet L=5e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.65e-07 covpccnr=0 wrxcnr=4.5e-06 sa=7.6e-07 sb=1.4e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M3@8 XI2/XI1/N1 XI2/N1N12 VSSA_RX VSSA_RX egnfet L=7e-07 W=9e-07
+ AD=6.3e-14 AS=6.3e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=8.1e-07 sa=9.6e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M2@3 XI2/XI1/VBP XI2/VBG XI2/XI1/N1 VSSA_RX egnfet L=5e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.65e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.4e-06 sb=7.6e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M3@7 XI2/XI1/N1 XI2/N1N12 VSSA_RX VSSA_RX egnfet L=7e-07 W=9e-07
+ AD=6.3e-14 AS=6.3e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=8.1e-07 sa=1.8e-06 sb=1.8e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M2@2 XI2/XI1/VBP XI2/VBG XI2/XI1/N1 VSSA_RX egnfet L=5e-07 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.65e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M3@6 XI2/XI1/N1 XI2/N1N12 VSSA_RX VSSA_RX egnfet L=7e-07 W=9e-07
+ AD=6.3e-14 AS=6.3e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06 sb=9.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M7 XI2/N1N12 XI2/N1N12 VSSA_RX VSSA_RX egnfet L=7e-07 W=9e-07
+ AD=1.08e-13 AS=6.3e-14 PD=2.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M1 XI2/XI1/N2 XI2/GMOUT XI2/XI1/N1 VSSA_RX egnfet L=5e-07 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.65e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M3@5 XI2/XI1/N1 XI2/N1N12 VSSA_RX VSSA_RX egnfet L=7e-07 W=9e-07
+ AD=6.3e-14 AS=1.08e-13 PD=1.04e-06 PS=2.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=8.1e-07 sa=1.2e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M1@4 XI2/XI1/N2 XI2/GMOUT XI2/XI1/N1 VSSA_RX egnfet L=5e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.65e-07 covpccnr=0 wrxcnr=4.5e-06 sa=7.6e-07 sb=1.4e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M3@4 XI2/XI1/N1 XI2/N1N12 VSSA_RX VSSA_RX egnfet L=7e-07 W=9e-07
+ AD=6.3e-14 AS=6.3e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=8.1e-07 sa=9.6e-07 sb=2.0083e-06 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M1@3 XI2/XI1/N2 XI2/GMOUT XI2/XI1/N1 VSSA_RX egnfet L=5e-07 W=5e-06
+ AD=3.5e-13 AS=3.5e-13 PD=5.14e-06 PS=5.14e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.65e-07 covpccnr=0 wrxcnr=4.5e-06 sa=1.4e-06 sb=7.6e-07 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M3@3 XI2/XI1/N1 XI2/N1N12 VSSA_RX VSSA_RX egnfet L=7e-07 W=9e-07
+ AD=6.3e-14 AS=6.3e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=8.1e-07 sa=1.8e-06 sb=1.8e-06 sd=0 ptwell=0
+ ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M1@2 XI2/XI1/N2 XI2/GMOUT XI2/XI1/N1 VSSA_RX egnfet L=5e-07 W=5e-06
+ AD=3.5e-13 AS=6e-13 PD=5.14e-06 PS=1.024e-05 M=1 sca=0 scb=0 scc=0
+ lpccnr=4.65e-07 covpccnr=0 wrxcnr=4.5e-06 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M3@2 XI2/XI1/N1 XI2/N1N12 VSSA_RX VSSA_RX egnfet L=7e-07 W=9e-07
+ AD=6.3e-14 AS=6.3e-14 PD=1.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06 sb=9.6e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M7@2 XI2/N1N12 XI2/N1N12 VSSA_RX VSSA_RX egnfet L=7e-07 W=9e-07
+ AD=1.08e-13 AS=6.3e-14 PD=2.04e-06 PS=1.04e-06 M=1 sca=0 scb=0 scc=0
+ lpccnr=6.45e-07 covpccnr=0 wrxcnr=8.1e-07 sa=2.0083e-06 sb=1.2e-07 sd=0
+ ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0 sizedup=0
+ pre_layout_local=0
XXI2/XI1/M13 VSSA_RX XI2/N1N12 VSSA_RX VSSA_RX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M13@4 VSSA_RX XI2/N1N12 VSSA_RX VSSA_RX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M13@3 VSSA_RX XI2/N1N12 VSSA_RX VSSA_RX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/M13@2 VSSA_RX XI2/N1N12 VSSA_RX VSSA_RX egnfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI2/XI1/XRR1/RR1 X290/X13/X7/noxref_6 XI2/GMOUT VDDHA_RX opppcres 2995.53 M=1
+ w=2e-06 l=9.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/XRR1/RR2 X290/X13/X7/noxref_6 X290/X13/X7/noxref_7 VDDHA_RX opppcres
+ 2995.53 M=1 w=2e-06 l=9.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/XRR1/RR3 X290/X13/X7/noxref_8 X290/X13/X7/noxref_7 VDDHA_RX opppcres
+ 2995.53 M=1 w=2e-06 l=9.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/XRR1/RR4 X290/X13/X7/noxref_8 X290/X13/X7/noxref_9 VDDHA_RX opppcres
+ 2995.53 M=1 w=2e-06 l=9.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/XRR1/RR5 X290/X13/X7/noxref_10 X290/X13/X7/noxref_9 VDDHA_RX opppcres
+ 2995.53 M=1 w=2e-06 l=9.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/XRR1/RR6 X290/X13/X7/noxref_10 X290/X13/X7/noxref_11 VDDHA_RX opppcres
+ 2995.53 M=1 w=2e-06 l=9.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/XRR1/RR7 X290/X13/X7/noxref_12 X290/X13/X7/noxref_11 VDDHA_RX opppcres
+ 2995.53 M=1 w=2e-06 l=9.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/XRR1/RR8 X290/X13/X7/noxref_12 X290/X13/X7/noxref_13 VDDHA_RX opppcres
+ 2995.53 M=1 w=2e-06 l=9.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/XRR1/RR9 X290/X13/X7/noxref_14 X290/X13/X7/noxref_13 VDDHA_RX opppcres
+ 2995.53 M=1 w=2e-06 l=9.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/XRR1/RR10 X290/X13/X7/noxref_14 VSSA_RX VDDHA_RX opppcres 2995.53 M=1
+ w=2e-06 l=9.8e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI1/MDC1@4 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@5 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@6 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@7 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@8 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@9 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@10 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@11 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=5.25548 scb=0.0046872
+ scc=0.000346407 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@12 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@13 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@14 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@15 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@16 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@17 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@18 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@19 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@20 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@21 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@22 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@23 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@24 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@25 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@26 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@27 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@28 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@29 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@30 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@31 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@32 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@33 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@34 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@35 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@36 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@37 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@38 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@39 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@40 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@41 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@42 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@43 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@44 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@45 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@46 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@47 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@48 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@49 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@50 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=0 scb=0 scc=0 lpccnr=4.515e-06
+ covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07 sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1
+ plorient=1 p_la=0 par=1 pccrit=0 sizedup=0 pre_layout_local=0
XXI1/MDC1@51 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=3.10078 scb=0.00278913
+ scc=0.000248935 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@52 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=5.25548 scb=0.0046872
+ scc=0.000346407 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@53 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@54 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@55 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@56 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@57 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@58 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=2.15471 scb=0.00189807
+ scc=9.74712e-05 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI1/MDC1@59 VDDHA_RX VSSA_RX VDDHA_RX VDDHA_RX egpfet L=5e-06 W=5e-06 AD=6e-13
+ AS=6e-13 PD=1.024e-05 PS=1.024e-05 M=1 sca=5.25548 scb=0.0046872
+ scc=0.000346407 lpccnr=4.515e-06 covpccnr=0 wrxcnr=4.5e-06 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=2 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI0/RRD1@2 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 5976.18 M=1 w=1e-06
+ l=9.72e-06   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI0/RRD1 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 5976.18 M=1 w=1e-06 l=9.72e-06
+ bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/RRD2@2 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 14482.7 M=1 w=1e-06
+ l=2.374e-05   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/RRD2 VDDHA_RX VDDHA_RX VDDHA_RX opppcres 14482.7 M=1 w=1e-06
+ l=2.374e-05   bp=1 pbar=1 s=1 ncr=1 sizedup=0
XXI2/XI1/CC0 XI2/GMOUT XI2/XI1/N1N209 VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC1 XI2/XI1/N1N209 XI2/GMOUT VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC2 XI2/GMOUT XI2/XI1/N1N209 VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC3 XI2/XI1/N1N209 XI2/GMOUT VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC4 XI2/GMOUT XI2/XI1/N1N209 VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC5 XI2/XI1/N1N209 XI2/GMOUT VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC6 XI2/GMOUT XI2/XI1/N1N209 VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC7 XI2/XI1/N1N209 XI2/GMOUT VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC8 XI2/GMOUT XI2/XI1/N1N209 VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC9 XI2/XI1/N1N209 XI2/GMOUT VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC10 XI2/GMOUT XI2/XI1/N1N209 VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC11 XI2/XI1/N1N209 XI2/GMOUT VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC12 XI2/GMOUT XI2/XI1/N1N209 VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/CC13 XI2/XI1/N1N209 XI2/GMOUT VSSA_RX vncap  botcap=0 botlev=17
+ setind=-2 toplev=31 sizedup=0 L=4.5e-06 W=3.78e-06
XXI2/XI1/X2I178/M0 XI2/XI1/X2I178/N1N42 XI2/XI1/X2I178/N1N42 VSSA_RX VSSA_RX
+ egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/X2I176/M0 XI2/XI1/X2I176/N1N42 XI2/XI1/X2I176/N1N42 VSSA_RX VSSA_RX
+ egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/X2I174/M0 XI2/XI1/X2I174/N1N42 XI2/XI1/X2I174/N1N42 VSSA_RX VSSA_RX
+ egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
XXI2/XI1/X2I171/M0 XI2/XI1/X2I171/N1N42 XI2/XI1/X2I171/N1N42 VSSA_RX VSSA_RX
+ egnfet L=1.5e-07 W=4e-07 AD=4.8e-14 AS=4.8e-14 PD=1.04e-06 PS=1.04e-06 M=1
+ sca=0 scb=0 scc=0 lpccnr=1.5e-07 covpccnr=0 wrxcnr=3.6e-07 sa=1.2e-07
+ sb=1.2e-07 sd=0 ptwell=0 ngcon=1 nf=1 plorient=1 p_la=0 par=1 pccrit=0
+ sizedup=0 pre_layout_local=0
c_141 VDD VSSA_RX:VSSA_TX:VSS 1.06419p
c_274 VSS VSSA_RX:VSSA_TX:VSS 1.08192p
c_455 VSSA_RX VSSA_RX:VSSA_TX:VSS 503.575f
c_607 VDDHA_RX VSSA_RX:VSSA_TX:VSS 390.515f
c_612 RXN VSSA_RX:VSSA_TX:VSS 8.10454f
c_617 RXP VSSA_RX:VSSA_TX:VSS 8.10127f
c_787 VDDHA_TX VSSA_RX:VSSA_TX:VSS 2.42066p
c_957 VSSA_TX VSSA_RX:VSSA_TX:VSS 1.76144p
c_968 TXP VSSA_RX:VSSA_TX:VSS 114.04f
c_979 TXN VSSA_RX:VSSA_TX:VSS 113.913f
c_999 PDRXI VSSA_RX:VSSA_TX:VSS 7.41902f
c_1014 DOI VSSA_RX:VSSA_TX:VSS 12.3545f
c_1045 IBRX2 VSSA_RX:VSSA_TX:VSS 11.7978f
c_1068 IBTX1 VSSA_RX:VSSA_TX:VSS 19.8327f
c_1080 CCMI0 VSSA_RX:VSSA_TX:VSS 2.48418f
c_1092 CCMI1 VSSA_RX:VSSA_TX:VSS 2.48418f
c_1104 CCMI2 VSSA_RX:VSSA_TX:VSS 2.48418f
c_1129 PDTXI VSSA_RX:VSSA_TX:VSS 7.05799f
c_1146 DTX VSSA_RX:VSSA_TX:VSS 1.12597f
c_1173 IBRX1 VSSA_RX:VSSA_TX:VSS 8.27098f
c_1183 CAI0 VSSA_RX:VSSA_TX:VSS 1.63915f
c_1193 CAI1 VSSA_RX:VSSA_TX:VSS 1.63915f
c_1203 CAI2 VSSA_RX:VSSA_TX:VSS 1.63915f
c_1222 PDI VSSA_RX:VSSA_TX:VSS 2.08494f
c_1326 IBTX2 VSSA_RX:VSSA_TX:VSS 30.4801f
c_1330 DO VSSA_RX:VSSA_TX:VSS 1.26612f
c_1336 CA0 VSSA_RX:VSSA_TX:VSS 0.994352f
c_1342 CA1 VSSA_RX:VSSA_TX:VSS 0.618821f
c_1348 CA2 VSSA_RX:VSSA_TX:VSS 0.613544f
c_1354 PD VSSA_RX:VSSA_TX:VSS 0.626462f
c_1360 PDTX VSSA_RX:VSSA_TX:VSS 0.640628f
c_1366 PDRX VSSA_RX:VSSA_TX:VSS 0.686397f
c_1372 CCM0 VSSA_RX:VSSA_TX:VSS 0.871795f
c_1378 CCM1 VSSA_RX:VSSA_TX:VSS 0.773638f
c_1384 CCM2 VSSA_RX:VSSA_TX:VSS 0.658814f
c_1392 LBEN VSSA_RX:VSSA_TX:VSS 0.772673f
c_1400 DI VSSA_RX:VSSA_TX:VSS 0.751255f
c_1415 XI1/VBP VSSA_RX:VSSA_TX:VSS 2.92197f
c_1433 XI1/INPI VSSA_RX:VSSA_TX:VSS 5.22338f
c_1451 XI1/INNI VSSA_RX:VSSA_TX:VSS 5.20992f
c_1463 XI1/INN1 VSSA_RX:VSSA_TX:VSS 1.91551f
c_1471 XI1/XI1/N0 VSSA_RX:VSSA_TX:VSS 0.869644f
c_1481 XI1/XI1/PDB VSSA_RX:VSSA_TX:VSS 1.00309f
c_1544 XI1/PDI VSSA_RX:VSSA_TX:VSS 9.02433f
c_1556 XI1/INP1 VSSA_RX:VSSA_TX:VSS 1.96615f
c_1570 XI1/XI5/O2 VSSA_RX:VSSA_TX:VSS 1.1331f
c_1583 XI1/XI5/O1 VSSA_RX:VSSA_TX:VSS 1.31214f
c_1589 XI1/XI3/X1I124/N1N50 VSSA_RX:VSSA_TX:VSS 0.155282f
c_1596 XI1/XI3/TIEL VSSA_RX:VSSA_TX:VSS 0.0956614f
c_1612 XI1/XI3/N2A VSSA_RX:VSSA_TX:VSS 0.63837f
c_1629 XI1/XI3/N2B VSSA_RX:VSSA_TX:VSS 0.647722f
c_1641 XI1/XI3/N1B VSSA_RX:VSSA_TX:VSS 0.56153f
c_1653 XI1/XI3/N1A VSSA_RX:VSSA_TX:VSS 0.567048f
c_1665 XI1/NN VSSA_RX:VSSA_TX:VSS 0.571999f
c_1673 XI1/XI3/N3B VSSA_RX:VSSA_TX:VSS 0.237244f
c_1685 XI1/NP VSSA_RX:VSSA_TX:VSS 0.58133f
c_1695 XI1/XI3/N3A VSSA_RX:VSSA_TX:VSS 0.373943f
c_1708 XI1/VAL VSSA_RX:VSSA_TX:VSS 1.13831f
c_1724 XI1/VBN VSSA_RX:VSSA_TX:VSS 1.7804f
c_1741 XI1/INP2 VSSA_RX:VSSA_TX:VSS 2.18331f
c_1758 XI1/INN2 VSSA_RX:VSSA_TX:VSS 1.93243f
c_1765 XI1/XI1/N1P VSSA_RX:VSSA_TX:VSS 0.71459f
c_1771 XI1/XI1/N2N VSSA_RX:VSSA_TX:VSS 0.472941f
c_1778 XI1/XI1/N1N VSSA_RX:VSSA_TX:VSS 0.71459f
c_1784 XI1/XI1/N2P VSSA_RX:VSSA_TX:VSS 0.472941f
c_1797 XI1/XI5/XI0B/PDB VSSA_RX:VSSA_TX:VSS 0.818508f
c_1807 XI1/XI5/XI0B/N1N422 VSSA_RX:VSSA_TX:VSS 0.400496f
c_1816 XI1/XI5/XI0B/N3P VSSA_RX:VSSA_TX:VSS 0.851582f
c_1825 XI1/XI5/XI0B/N3N VSSA_RX:VSSA_TX:VSS 0.855316f
c_1833 XI1/XI5/XI0B/N0 VSSA_RX:VSSA_TX:VSS 0.691052f
c_1841 XI1/XI5/XI0B/N2P VSSA_RX:VSSA_TX:VSS 0.324078f
c_1850 XI1/XI5/XI0B/N1N VSSA_RX:VSSA_TX:VSS 0.536655f
c_1859 XI1/XI5/XI0B/N2N VSSA_RX:VSSA_TX:VSS 0.329663f
c_1868 XI1/XI5/XI0B/N1P VSSA_RX:VSSA_TX:VSS 0.537417f
c_1881 XI1/XI5/XI0A/PDB VSSA_RX:VSSA_TX:VSS 0.819718f
c_1891 XI1/XI5/XI0A/N1N422 VSSA_RX:VSSA_TX:VSS 0.400496f
c_1900 XI1/XI5/XI0A/N3P VSSA_RX:VSSA_TX:VSS 0.851609f
c_1909 XI1/XI5/XI0A/N3N VSSA_RX:VSSA_TX:VSS 0.855316f
c_1917 XI1/XI5/XI0A/N0 VSSA_RX:VSSA_TX:VSS 0.51549f
c_1925 XI1/XI5/XI0A/N2P VSSA_RX:VSSA_TX:VSS 0.324086f
c_1934 XI1/XI5/XI0A/N1N VSSA_RX:VSSA_TX:VSS 0.551173f
c_1943 XI1/XI5/XI0A/N2N VSSA_RX:VSSA_TX:VSS 0.329671f
c_1951 XI1/XI5/XI0A/N1P VSSA_RX:VSSA_TX:VSS 0.551952f
c_1956 XI1/XI3/XG3B/N1 VSSA_RX:VSSA_TX:VSS 3.00226e-19
c_1962 XI1/XI3/XG3A/N1 VSSA_RX:VSSA_TX:VSS 5.01334e-19
c_1970 XI1/XI3/N4A VSSA_RX:VSSA_TX:VSS 0.475547f
c_1978 XI1/XI3/N5A VSSA_RX:VSSA_TX:VSS 0.704841f
c_1984 XI1/XI5/N1N356 VSSA_RX:VSSA_TX:VSS 0.306569f
c_1989 XI1/XI5/XG0/N1 VSSA_RX:VSSA_TX:VSS 7.71098e-19
c_1997 XI1/XI5/N1N284 VSSA_RX:VSSA_TX:VSS 0.287016f
c_2001 XI1/XI5/N1N312 VSSA_RX:VSSA_TX:VSS 0.435254f
c_2006 X286/X88/noxref_55 VSSA_RX:VSSA_TX:VSS 0.194079f
c_2011 X286/X88/noxref_56 VSSA_RX:VSSA_TX:VSS 0.195095f
c_2015 X286/X88/noxref_57 VSSA_RX:VSSA_TX:VSS 0.219277f
c_2035 XI1/XI4/PDB VSSA_RX:VSSA_TX:VSS 1.07769f
c_2048 XI1/XI4/N1N VSSA_RX:VSSA_TX:VSS 0.349039f
c_2061 XI1/XI4/N1P VSSA_RX:VSSA_TX:VSS 0.369688f
c_2067 XI1/XI6/N1N36 VSSA_RX:VSSA_TX:VSS 0.360094f
c_2075 XI1/XI6/N1N5 VSSA_RX:VSSA_TX:VSS 0.36317f
c_2083 XI1/XI6/N2 VSSA_RX:VSSA_TX:VSS 0.518289f
c_2091 XI1/XI6/N1 VSSA_RX:VSSA_TX:VSS 0.452363f
c_2097 XI1/XI6/N3 VSSA_RX:VSSA_TX:VSS 1.09571f
c_2108 XI1/XI2/PDIB VSSA_RX:VSSA_TX:VSS 1.27619f
c_2120 XI1/XI2/PDI VSSA_RX:VSSA_TX:VSS 0.994478f
c_2130 XI1/XI2/N1N204 VSSA_RX:VSSA_TX:VSS 1.2237f
c_2140 XI1/XI2/N1N VSSA_RX:VSSA_TX:VSS 0.75871f
c_2150 XI1/XI2/N1P VSSA_RX:VSSA_TX:VSS 0.758896f
c_2162 XI1/XI0/N7 VSSA_RX:VSSA_TX:VSS 1.41245f
c_2170 XI1/XI0/PDB VSSA_RX:VSSA_TX:VSS 0.339794f
c_2174 XI1/XI0/N3 VSSA_RX:VSSA_TX:VSS 0.0539459f
c_2187 XI1/XI0/N2 VSSA_RX:VSSA_TX:VSS 1.51835f
c_2192 XI1/XI0/N4 VSSA_RX:VSSA_TX:VSS 0.0256126f
c_2197 XI1/XI0/N8 VSSA_RX:VSSA_TX:VSS 0.0495098f
c_2203 XI1/XI0/N6 VSSA_RX:VSSA_TX:VSS 0.039523f
c_2209 XI1/XI0/N9 VSSA_RX:VSSA_TX:VSS 0.0275825f
c_2215 XI1/XI0/N10 VSSA_RX:VSSA_TX:VSS 0.0206592f
c_2254 XI0/CCMH0 VSSA_RX:VSSA_TX:VSS 3.79524f
c_2289 XI0/CCMH1 VSSA_RX:VSSA_TX:VSS 4.20159f
c_2297 XI0/PDH VSSA_RX:VSSA_TX:VSS 3.78866f
c_2325 XI0/EN VSSA_RX:VSSA_TX:VSS 2.60062f
c_2362 XI0/CCMH2 VSSA_RX:VSSA_TX:VSS 5.29995f
c_2388 XI0/VBP VSSA_RX:VSSA_TX:VSS 171.966f
c_2447 XI0/VCM VSSA_RX:VSSA_TX:VSS 43.1397f
c_2458 XI0/XI1/N1N166 VSSA_RX:VSSA_TX:VSS 88.7029f
c_2482 XI0/FB VSSA_RX:VSSA_TX:VSS 1.93103f
c_2494 XI0/XI1/XI0/VCM7 VSSA_RX:VSSA_TX:VSS 0.489738f
c_2511 XI0/XI1/XI0/VCM6 VSSA_RX:VSSA_TX:VSS 0.666357f
c_2527 XI0/XI1/XI0/VCM5 VSSA_RX:VSSA_TX:VSS 0.492414f
c_2544 XI0/XI1/XI0/VCM4 VSSA_RX:VSSA_TX:VSS 0.761041f
c_2557 XI0/XI1/XI0/VCM3 VSSA_RX:VSSA_TX:VSS 0.493904f
c_2572 XI0/XI1/XI0/VCM2 VSSA_RX:VSSA_TX:VSS 0.705881f
c_2585 XI0/XI1/XI0/VCM1 VSSA_RX:VSSA_TX:VSS 0.493277f
c_2598 XI0/XI1/XI0/VCM0 VSSA_RX:VSSA_TX:VSS 1.124f
c_2617 XI0/XI1/XI1/N6 VSSA_RX:VSSA_TX:VSS 2.25962f
c_2638 XI0/XI1/PD VSSA_RX:VSSA_TX:VSS 1.50624f
c_2651 XI0/XI1/XI1/N7 VSSA_RX:VSSA_TX:VSS 1.26501f
c_2663 XI0/XI1/XI1/N14 VSSA_RX:VSSA_TX:VSS 1.29281f
c_2680 XI0/XI1/XI1/N10 VSSA_RX:VSSA_TX:VSS 1.13595f
c_2689 XI0/XI1/XI1/N3 VSSA_RX:VSSA_TX:VSS 0.262297f
c_2709 XI0/XI1/XI1/N9 VSSA_RX:VSSA_TX:VSS 1.41708f
c_2725 XI0/XI1/XI1/N8 VSSA_RX:VSSA_TX:VSS 1.87696f
c_2733 XI0/XI1/N1N69 VSSA_RX:VSSA_TX:VSS 0.380078f
c_2735 X287/X22/X117/noxref_11 VSSA_RX:VSSA_TX:VSS 0.216284f
c_2740 XI0/XI1/N1 VSSA_RX:VSSA_TX:VSS 0.546091f
c_2744 X287/X22/X118/noxref_13 VSSA_RX:VSSA_TX:VSS 0.231266f
c_2749 X287/X22/X118/noxref_14 VSSA_RX:VSSA_TX:VSS 0.0413205f
c_2753 X287/X22/X118/noxref_15 VSSA_RX:VSSA_TX:VSS 0.232478f
c_2758 X287/X22/X118/noxref_16 VSSA_RX:VSSA_TX:VSS 0.0432745f
c_2762 X287/X22/X118/noxref_17 VSSA_RX:VSSA_TX:VSS 0.233559f
c_2767 X287/X22/X118/noxref_18 VSSA_RX:VSSA_TX:VSS 0.0413047f
c_2770 X287/X22/X118/noxref_19 VSSA_RX:VSSA_TX:VSS 0.231393f
c_2777 XI0/XI1/XI0/XI0/N1N140 VSSA_RX:VSSA_TX:VSS 0.373403f
c_2785 XI0/XI1/XI0/XI0/N1N134 VSSA_RX:VSSA_TX:VSS 0.367774f
c_2814 XI0/XI1/XI0/XI0/COI VSSA_RX:VSSA_TX:VSS 2.30246f
c_2842 XI0/XI1/XI0/XI0/C1I VSSA_RX:VSSA_TX:VSS 2.35194f
c_2865 XI0/XI1/XI0/XI0/SHB VSSA_RX:VSSA_TX:VSS 0.467685f
c_2887 XI0/XI1/XI0/XI0/SH VSSA_RX:VSSA_TX:VSS 0.379158f
c_2906 XI0/XI1/XI0/XI0/N1 VSSA_RX:VSSA_TX:VSS 0.449959f
c_2916 XI0/XI1/XI0/XI0/XI1/C0B VSSA_RX:VSSA_TX:VSS 0.339612f
c_2936 XI0/XI1/XI0/XI0/XI1/S3 VSSA_RX:VSSA_TX:VSS 0.651543f
c_2946 XI0/XI1/XI0/XI0/XI1/C1B VSSA_RX:VSSA_TX:VSS 0.369474f
c_2967 XI0/XI1/XI0/XI0/XI1/S2 VSSA_RX:VSSA_TX:VSS 0.615979f
c_2988 XI0/XI1/XI0/XI0/XI1/S1 VSSA_RX:VSSA_TX:VSS 0.580421f
c_2999 XI0/XI1/XI0/XI0/XI1/S0 VSSA_RX:VSSA_TX:VSS 0.122022f
c_3010 XI0/XI1/XI0/XI0/XI1/N1 VSSA_RX:VSSA_TX:VSS 0.325752f
c_3028 XI0/XI1/XI0/XI0/XI1/S0B VSSA_RX:VSSA_TX:VSS 0.628539f
c_3039 XI0/XI1/XI0/XI0/XI1/S3B VSSA_RX:VSSA_TX:VSS 0.0870004f
c_3051 XI0/XI1/XI0/XI0/XI1/S2B VSSA_RX:VSSA_TX:VSS 0.0869697f
c_3063 XI0/XI1/XI0/XI0/XI1/S1B VSSA_RX:VSSA_TX:VSS 0.0869697f
c_3073 XI0/XI1/XI0/XI0/XI1/N4 VSSA_RX:VSSA_TX:VSS 0.326002f
c_3084 XI0/XI1/XI0/XI0/XI1/N3 VSSA_RX:VSSA_TX:VSS 0.328036f
c_3095 XI0/XI1/XI0/XI0/XI1/N2 VSSA_RX:VSSA_TX:VSS 0.327025f
c_3124 XI0/XI1/XI0/XI0/N2 VSSA_RX:VSSA_TX:VSS 0.473891f
c_3134 XI0/XI1/XI0/XI0/XI0/C0B VSSA_RX:VSSA_TX:VSS 0.339612f
c_3153 XI0/XI1/XI0/XI0/XI0/S3 VSSA_RX:VSSA_TX:VSS 0.652485f
c_3163 XI0/XI1/XI0/XI0/XI0/C1B VSSA_RX:VSSA_TX:VSS 0.369474f
c_3182 XI0/XI1/XI0/XI0/XI0/S2 VSSA_RX:VSSA_TX:VSS 0.616921f
c_3201 XI0/XI1/XI0/XI0/XI0/S1 VSSA_RX:VSSA_TX:VSS 0.581363f
c_3210 XI0/XI1/XI0/XI0/XI0/S0 VSSA_RX:VSSA_TX:VSS 0.122817f
c_3221 XI0/XI1/XI0/XI0/XI0/N1 VSSA_RX:VSSA_TX:VSS 0.325232f
c_3236 XI0/XI1/XI0/XI0/XI0/S0B VSSA_RX:VSSA_TX:VSS 0.675194f
c_3246 XI0/XI1/XI0/XI0/XI0/S3B VSSA_RX:VSSA_TX:VSS 0.0877953f
c_3256 XI0/XI1/XI0/XI0/XI0/S2B VSSA_RX:VSSA_TX:VSS 0.0877646f
c_3266 XI0/XI1/XI0/XI0/XI0/S1B VSSA_RX:VSSA_TX:VSS 0.0877646f
c_3277 XI0/XI1/XI0/XI0/XI0/N4 VSSA_RX:VSSA_TX:VSS 0.32779f
c_3288 XI0/XI1/XI0/XI0/XI0/N3 VSSA_RX:VSSA_TX:VSS 0.328036f
c_3299 XI0/XI1/XI0/XI0/XI0/N2 VSSA_RX:VSSA_TX:VSS 0.327025f
c_3319 XI0/XI1/XI1/XI0/N4 VSSA_RX:VSSA_TX:VSS 0.280999f
c_3326 XI0/XI1/XI1/XI0/N1N5 VSSA_RX:VSSA_TX:VSS 0.0303487f
c_3338 XI0/XI1/XI1/XI0/N2 VSSA_RX:VSSA_TX:VSS 0.678871f
c_3349 XI0/XI1/XI1/XI0/TIEL VSSA_RX:VSSA_TX:VSS 0.241099f
c_3358 XI0/XI1/XI1/XI0/X1I44/N1N50 VSSA_RX:VSSA_TX:VSS 0.167872f
c_3364 XI0/XI1/XI1/XI0/N3 VSSA_RX:VSSA_TX:VSS 0.469501f
c_3368 XI0/XI1/XI1/N1N21 VSSA_RX:VSSA_TX:VSS 0.0481451f
c_3373 XI0/XI1/XI1/N1N4 VSSA_RX:VSSA_TX:VSS 0.0373142f
c_3376 XI0/XI1/XI1/N1N22 VSSA_RX:VSSA_TX:VSS 0.039085f
c_3380 XI0/XI1/XI1/N1N24 VSSA_RX:VSSA_TX:VSS 0.0524008f
c_3384 XI0/XI1/XI1/N4 VSSA_RX:VSSA_TX:VSS 0.246684f
c_3397 XI0/XI1/XI1/N1 VSSA_RX:VSSA_TX:VSS 0.434274f
c_3402 XI0/XI1/XI1/N5 VSSA_RX:VSSA_TX:VSS 0.246684f
c_3415 XI0/XI1/XI1/N2 VSSA_RX:VSSA_TX:VSS 0.439354f
c_3424 XI0/XI1/PDB VSSA_RX:VSSA_TX:VSS 0.298886f
c_3429 XI0/N1N229 VSSA_RX:VSSA_TX:VSS 0.217164f
c_3439 XI0/N1N225 VSSA_RX:VSSA_TX:VSS 1.0091f
c_3444 XI0/XI3A0/N1N36 VSSA_RX:VSSA_TX:VSS 0.304461f
c_3450 XI0/XI3A0/N1N5 VSSA_RX:VSSA_TX:VSS 0.279601f
c_3457 XI0/XI3A0/N2 VSSA_RX:VSSA_TX:VSS 0.465359f
c_3464 XI0/XI3A0/N1 VSSA_RX:VSSA_TX:VSS 0.404749f
c_3472 XI0/XI3A0/N3 VSSA_RX:VSSA_TX:VSS 0.558857f
c_3477 XI0/XI3A1/N1N36 VSSA_RX:VSSA_TX:VSS 0.304461f
c_3483 XI0/XI3A1/N1N5 VSSA_RX:VSSA_TX:VSS 0.279601f
c_3490 XI0/XI3A1/N2 VSSA_RX:VSSA_TX:VSS 0.465359f
c_3497 XI0/XI3A1/N1 VSSA_RX:VSSA_TX:VSS 0.404749f
c_3505 XI0/XI3A1/N3 VSSA_RX:VSSA_TX:VSS 0.558857f
c_3510 XI0/XI3A2/N1N36 VSSA_RX:VSSA_TX:VSS 0.304461f
c_3516 XI0/XI3A2/N1N5 VSSA_RX:VSSA_TX:VSS 0.279601f
c_3523 XI0/XI3A2/N2 VSSA_RX:VSSA_TX:VSS 0.465359f
c_3530 XI0/XI3A2/N1 VSSA_RX:VSSA_TX:VSS 0.404749f
c_3538 XI0/XI3A2/N3 VSSA_RX:VSSA_TX:VSS 0.558857f
c_3543 XI0/XI2/N1N36 VSSA_RX:VSSA_TX:VSS 0.304461f
c_3549 XI0/XI2/N1N5 VSSA_RX:VSSA_TX:VSS 0.279601f
c_3556 XI0/XI2/N2 VSSA_RX:VSSA_TX:VSS 0.465359f
c_3563 XI0/XI2/N1 VSSA_RX:VSSA_TX:VSS 0.404749f
c_3572 XI0/XI2/N3 VSSA_RX:VSSA_TX:VSS 0.526459f
c_3581 XI0/XI0/XI2/PDB VSSA_RX:VSSA_TX:VSS 0.915311f
c_3607 XI0/XI0/ENBH VSSA_RX:VSSA_TX:VSS 7.71284f
c_3620 XI0/XI0/NN3B VSSA_RX:VSSA_TX:VSS 24.4343f
c_3633 XI0/XI0/NN3A VSSA_RX:VSSA_TX:VSS 23.2044f
c_3646 XI0/XI0/NP3A VSSA_RX:VSSA_TX:VSS 21.0652f
c_3659 XI0/XI0/NP3B VSSA_RX:VSSA_TX:VSS 22.6017f
c_3674 XI0/XI0/NP1 VSSA_RX:VSSA_TX:VSS 0.980014f
c_3689 XI0/XI0/NN1 VSSA_RX:VSSA_TX:VSS 0.9244f
c_3701 XI0/XI0/NP2 VSSA_RX:VSSA_TX:VSS 0.637834f
c_3713 XI0/XI0/NN2 VSSA_RX:VSSA_TX:VSS 0.637672f
c_3718 XI0/XI0/XI2/X1I43/N1N36 VSSA_RX:VSSA_TX:VSS 0.309433f
c_3724 XI0/XI0/XI2/X1I43/N1N5 VSSA_RX:VSSA_TX:VSS 0.280756f
c_3731 XI0/XI0/XI2/X1I43/N2 VSSA_RX:VSSA_TX:VSS 0.471107f
c_3738 XI0/XI0/XI2/X1I43/N1 VSSA_RX:VSSA_TX:VSS 0.410612f
c_3746 XI0/XI0/XI2/X1I43/N3 VSSA_RX:VSSA_TX:VSS 0.560517f
c_3763 XI0/XI0/XI3/TIEH VSSA_RX:VSSA_TX:VSS 0.393491f
c_3769 XI0/XI0/XI3/X1I221/N1N42 VSSA_RX:VSSA_TX:VSS 0.181603f
c_3780 XI0/XI0/XI3/N0N VSSA_RX:VSSA_TX:VSS 1.00664f
c_3793 XI0/XI0/XI3/TIEL VSSA_RX:VSSA_TX:VSS 0.232261f
c_3804 XI0/XI0/XI3/N0P VSSA_RX:VSSA_TX:VSS 0.904052f
c_3811 XI0/XI0/XI3/X1I218/N1N50 VSSA_RX:VSSA_TX:VSS 0.135799f
c_3820 XI0/XI0/XI3/NN VSSA_RX:VSSA_TX:VSS 0.715397f
c_3830 XI0/XI0/XI3/NP VSSA_RX:VSSA_TX:VSS 0.658301f
c_3840 XI0/XI0/XI3/N1N206 VSSA_RX:VSSA_TX:VSS 0.467929f
c_3852 XI0/XI0/XI3/N1N207 VSSA_RX:VSSA_TX:VSS 0.407804f
c_3867 XI0/XI0/XI3/IN4 VSSA_RX:VSSA_TX:VSS 0.823493f
c_3876 XI0/XI0/XI3/IN1 VSSA_RX:VSSA_TX:VSS 0.210893f
c_3884 XI0/XI0/XI3/IN2 VSSA_RX:VSSA_TX:VSS 0.246328f
c_3891 XI0/XI0/XI3/IN3 VSSA_RX:VSSA_TX:VSS 0.392553f
c_3902 XI0/XI0/XI2/N1 VSSA_RX:VSSA_TX:VSS 0.305627f
c_3910 XI0/XI0/XI2/N2 VSSA_RX:VSSA_TX:VSS 0.300799f
c_3932 XI0/XI0/CM VSSA_RX:VSSA_TX:VSS 107.463f
c_3940 XI0/XI0/XI0/XI0/N1N152 VSSA_RX:VSSA_TX:VSS 1.14546f
c_3949 XI0/XI0/XI0/XI0/N2N VSSA_RX:VSSA_TX:VSS 0.420254f
c_3966 XI0/XI0/XI0/VBN VSSA_RX:VSSA_TX:VSS 14.4274f
c_3972 XI0/XI0/XI0/N3 VSSA_RX:VSSA_TX:VSS 83.1684f
c_3981 XI0/XI0/XI0/XI0/N1 VSSA_RX:VSSA_TX:VSS 3.04061f
c_3993 XI0/XI0/XI0/N2 VSSA_RX:VSSA_TX:VSS 72.9012f
c_4008 XI0/XI0/XI0/N1 VSSA_RX:VSSA_TX:VSS 116.682f
c_4013 XI0/XI0/XI0/N1N798 VSSA_RX:VSSA_TX:VSS 0.0422157f
c_4018 XI0/XI0/XI0/N1N789 VSSA_RX:VSSA_TX:VSS 0.0358448f
c_4024 XI0/XI0/XI1/N1N118 VSSA_RX:VSSA_TX:VSS 0.225795f
c_4060 XI0/XI0/XI1/S1B VSSA_RX:VSSA_TX:VSS 3.01929f
c_4096 XI0/XI0/XI1/S1 VSSA_RX:VSSA_TX:VSS 2.80852f
c_4102 XI0/XI0/XI1/NN VSSA_RX:VSSA_TX:VSS 0.26112f
c_4109 XI0/XI0/XI1/NP VSSA_RX:VSSA_TX:VSS 0.444104f
c_4126 XI0/XI0/XI1/N1 VSSA_RX:VSSA_TX:VSS 1.31031f
c_4137 XI0/XI0/XI1/XI1P/N1N29 VSSA_RX:VSSA_TX:VSS 0.171896f
c_4145 XI0/XI0/XI1/XI1P/N1N28 VSSA_RX:VSSA_TX:VSS 0.430161f
c_4153 XI0/XI0/XI1/XI1P/N1N25 VSSA_RX:VSSA_TX:VSS 0.703602f
c_4159 XI0/XI0/XI1/XI1P/N1N42 VSSA_RX:VSSA_TX:VSS 6.05103e-19
c_4163 XI0/XI0/XI1/XI1P/N1N50 VSSA_RX:VSSA_TX:VSS 7.93718e-19
c_4169 XI0/XI0/XI1/XI1P/N1N38 VSSA_RX:VSSA_TX:VSS 0.00207689f
c_4174 XI0/XI0/XI1/XI1P/N1N52 VSSA_RX:VSSA_TX:VSS 0.00230825f
c_4185 XI0/XI0/XI1/XI0P/N1N29 VSSA_RX:VSSA_TX:VSS 0.164309f
c_4193 XI0/XI0/XI1/XI0P/N1N28 VSSA_RX:VSSA_TX:VSS 0.415884f
c_4201 XI0/XI0/XI1/XI0P/N1N25 VSSA_RX:VSSA_TX:VSS 0.727816f
c_4207 XI0/XI0/XI1/XI0P/N1N42 VSSA_RX:VSSA_TX:VSS 6.05103e-19
c_4212 XI0/XI0/XI1/XI0P/N1N50 VSSA_RX:VSSA_TX:VSS 7.93718e-19
c_4218 XI0/XI0/XI1/XI0P/N1N38 VSSA_RX:VSSA_TX:VSS 6.85616e-19
c_4222 XI0/XI0/XI1/XI0P/N1N52 VSSA_RX:VSSA_TX:VSS 0.00315511f
c_4239 XI0/XI0/XI1/N2 VSSA_RX:VSSA_TX:VSS 1.32074f
c_4250 XI0/XI0/XI1/XI1N/N1N29 VSSA_RX:VSSA_TX:VSS 0.173237f
c_4258 XI0/XI0/XI1/XI1N/N1N28 VSSA_RX:VSSA_TX:VSS 0.432345f
c_4266 XI0/XI0/XI1/XI1N/N1N25 VSSA_RX:VSSA_TX:VSS 0.710267f
c_4272 XI0/XI0/XI1/XI1N/N1N42 VSSA_RX:VSSA_TX:VSS 6.05103e-19
c_4276 XI0/XI0/XI1/XI1N/N1N50 VSSA_RX:VSSA_TX:VSS 7.93718e-19
c_4282 XI0/XI0/XI1/XI1N/N1N38 VSSA_RX:VSSA_TX:VSS 0.00292375f
c_4287 XI0/XI0/XI1/XI1N/N1N52 VSSA_RX:VSSA_TX:VSS 0.00315511f
c_4298 XI0/XI0/XI1/XI0N/N1N29 VSSA_RX:VSSA_TX:VSS 0.165001f
c_4306 XI0/XI0/XI1/XI0N/N1N28 VSSA_RX:VSSA_TX:VSS 0.416576f
c_4314 XI0/XI0/XI1/XI0N/N1N25 VSSA_RX:VSSA_TX:VSS 0.729892f
c_4320 XI0/XI0/XI1/XI0N/N1N42 VSSA_RX:VSSA_TX:VSS 6.05103e-19
c_4325 XI0/XI0/XI1/XI0N/N1N50 VSSA_RX:VSSA_TX:VSS 7.93718e-19
c_4331 XI0/XI0/XI1/XI0N/N1N38 VSSA_RX:VSSA_TX:VSS 6.85616e-19
c_4335 XI0/XI0/XI1/XI0N/N1N52 VSSA_RX:VSSA_TX:VSS 0.00315511f
c_4371 DLBI VSSA_RX:VSSA_TX:VSS 3.45726f
c_4390 DLB VSSA_RX:VSSA_TX:VSS 3.26083f
c_4402 N1N291 VSSA_RX:VSSA_TX:VSS 0.338963f
c_4409 XI3/N1 VSSA_RX:VSSA_TX:VSS 0.190884f
c_4417 XI4/SLB VSSA_RX:VSSA_TX:VSS 0.249321f
c_4427 XI4/SL VSSA_RX:VSSA_TX:VSS 0.191163f
c_4437 XI4/N1 VSSA_RX:VSSA_TX:VSS 0.17518f
c_4445 XI4/N2 VSSA_RX:VSSA_TX:VSS 0.143421f
c_4456 XI9A0/N2 VSSA_RX:VSSA_TX:VSS 0.230587f
c_4462 XI9A1/N2 VSSA_RX:VSSA_TX:VSS 0.230587f
c_4468 XI9A2/N2 VSSA_RX:VSSA_TX:VSS 0.230587f
c_4474 XI8/N2 VSSA_RX:VSSA_TX:VSS 0.230053f
c_4480 XI5A0/N2 VSSA_RX:VSSA_TX:VSS 0.230587f
c_4486 XI5A1/N2 VSSA_RX:VSSA_TX:VSS 0.230587f
c_4492 XI5A2/N2 VSSA_RX:VSSA_TX:VSS 0.230587f
c_4499 XI12/N2 VSSA_RX:VSSA_TX:VSS 0.228272f
c_4506 XI12/N3 VSSA_RX:VSSA_TX:VSS 0.518685f
c_4511 XI12/N4 VSSA_RX:VSSA_TX:VSS 0.655383f
c_4517 XI11/N2 VSSA_RX:VSSA_TX:VSS 0.230146f
c_4525 XI11/N3 VSSA_RX:VSSA_TX:VSS 0.518108f
c_4531 XI11/N4 VSSA_RX:VSSA_TX:VSS 0.655f
c_4542 XI6/N0 VSSA_RX:VSSA_TX:VSS 0.177957f
c_4550 XI6/N1 VSSA_RX:VSSA_TX:VSS 0.18257f
c_4559 XI6/N2 VSSA_RX:VSSA_TX:VSS 0.227698f
c_4568 XI6/N3 VSSA_RX:VSSA_TX:VSS 0.514984f
c_4575 XI6/N4 VSSA_RX:VSSA_TX:VSS 0.645578f
c_4587 XI7/N0 VSSA_RX:VSSA_TX:VSS 0.178671f
c_4594 XI7/N1 VSSA_RX:VSSA_TX:VSS 0.184031f
c_4602 XI7/N2 VSSA_RX:VSSA_TX:VSS 0.229123f
c_4611 XI7/N3 VSSA_RX:VSSA_TX:VSS 0.515713f
c_4618 XI7/N4 VSSA_RX:VSSA_TX:VSS 0.647138f
c_4625 XI10/N2 VSSA_RX:VSSA_TX:VSS 0.227953f
c_4631 XI10/N3 VSSA_RX:VSSA_TX:VSS 0.518271f
c_4636 XI10/N4 VSSA_RX:VSSA_TX:VSS 0.652204f
c_4678 XI2/PDI VSSA_RX:VSSA_TX:VSS 3.69494f
c_4707 XI2/PDTXI VSSA_RX:VSSA_TX:VSS 2.66844f
c_4725 XI2/PDRXI VSSA_RX:VSSA_TX:VSS 1.7119f
c_4757 XI2/CAI2 VSSA_RX:VSSA_TX:VSS 1.80318f
c_4789 XI2/CAI1 VSSA_RX:VSSA_TX:VSS 1.70041f
c_4802 XI2/N1N12 VSSA_RX:VSSA_TX:VSS 2.66137f
c_4834 XI2/CAI0 VSSA_RX:VSSA_TX:VSS 1.75379f
c_4857 XI2/VBG VSSA_RX:VSSA_TX:VSS 3.04293f
c_4863 XI2/XI3/N1N36 VSSA_RX:VSSA_TX:VSS 0.483293f
c_4870 XI2/XI3/N1N5 VSSA_RX:VSSA_TX:VSS 0.539529f
c_4877 XI2/XI3/N2 VSSA_RX:VSSA_TX:VSS 0.627565f
c_4884 XI2/XI3/N1 VSSA_RX:VSSA_TX:VSS 0.610195f
c_4891 XI2/XI3/N3 VSSA_RX:VSSA_TX:VSS 0.443988f
c_4897 XI2/XI4/N1N36 VSSA_RX:VSSA_TX:VSS 0.483428f
c_4904 XI2/XI4/N1N5 VSSA_RX:VSSA_TX:VSS 0.539529f
c_4911 XI2/XI4/N2 VSSA_RX:VSSA_TX:VSS 0.627565f
c_4918 XI2/XI4/N1 VSSA_RX:VSSA_TX:VSS 0.610195f
c_4925 XI2/XI4/N3 VSSA_RX:VSSA_TX:VSS 0.447224f
c_4931 XI2/XI2/N1N36 VSSA_RX:VSSA_TX:VSS 0.483399f
c_4938 XI2/XI2/N1N5 VSSA_RX:VSSA_TX:VSS 0.539529f
c_4945 XI2/XI2/N2 VSSA_RX:VSSA_TX:VSS 0.627565f
c_4952 XI2/XI2/N1 VSSA_RX:VSSA_TX:VSS 0.610195f
c_4959 XI2/XI2/N3 VSSA_RX:VSSA_TX:VSS 0.447224f
c_4965 XI2/XI5A2/N1N36 VSSA_RX:VSSA_TX:VSS 0.486822f
c_4972 XI2/XI5A2/N1N5 VSSA_RX:VSSA_TX:VSS 0.539529f
c_4979 XI2/XI5A2/N2 VSSA_RX:VSSA_TX:VSS 0.627565f
c_4986 XI2/XI5A2/N1 VSSA_RX:VSSA_TX:VSS 0.610195f
c_4993 XI2/XI5A2/N3 VSSA_RX:VSSA_TX:VSS 0.447224f
c_5000 XI2/XI5A1/N1N36 VSSA_RX:VSSA_TX:VSS 0.485473f
c_5008 XI2/XI5A1/N1N5 VSSA_RX:VSSA_TX:VSS 0.536534f
c_5016 XI2/XI5A1/N2 VSSA_RX:VSSA_TX:VSS 0.62527f
c_5024 XI2/XI5A1/N1 VSSA_RX:VSSA_TX:VSS 0.607274f
c_5031 XI2/XI5A1/N3 VSSA_RX:VSSA_TX:VSS 0.447224f
c_5039 XI2/XI5A0/N1N36 VSSA_RX:VSSA_TX:VSS 0.484167f
c_5048 XI2/XI5A0/N1N5 VSSA_RX:VSSA_TX:VSS 0.533539f
c_5057 XI2/XI5A0/N2 VSSA_RX:VSSA_TX:VSS 0.622975f
c_5066 XI2/XI5A0/N1 VSSA_RX:VSSA_TX:VSS 0.604353f
c_5073 XI2/XI5A0/N3 VSSA_RX:VSSA_TX:VSS 0.447224f
c_5088 XI2/XI0/INP VSSA_RX:VSSA_TX:VSS 0.91629f
c_5095 XI2/XI0/N1 VSSA_RX:VSSA_TX:VSS 9.02355f
c_5102 XI2/XI0/N2 VSSA_RX:VSSA_TX:VSS 5.76978f
c_5119 XI2/XI0/INN VSSA_RX:VSSA_TX:VSS 1.91337f
c_5145 XI2/VBP VSSA_RX:VSSA_TX:VSS 8.28983f
c_5161 XI2/XI0/XOP/N6 VSSA_RX:VSSA_TX:VSS 3.18474f
c_5176 XI2/XI0/XOP/N14 VSSA_RX:VSSA_TX:VSS 1.54223f
c_5186 XI2/XI0/PDB VSSA_RX:VSSA_TX:VSS 0.634525f
c_5195 XI2/XI0/N3 VSSA_RX:VSSA_TX:VSS 0.145235f
c_5200 XI2/XI0/XG2/N1 VSSA_RX:VSSA_TX:VSS 0.00731482f
c_5204 X290/X12/X50/noxref_8 VSSA_RX:VSSA_TX:VSS 0.0349658f
c_5206 X290/X12/X50/noxref_9 VSSA_RX:VSSA_TX:VSS 0.0363402f
c_5210 X290/X12/X50/X4/noxref_5 VSSA_RX:VSSA_TX:VSS 0.0922163f
c_5214 X290/X12/X50/X4/noxref_6 VSSA_RX:VSSA_TX:VSS 0.115606f
c_5219 X290/X12/X50/X4/noxref_7 VSSA_RX:VSSA_TX:VSS 0.0929123f
c_5222 X290/X12/X50/X4/noxref_8 VSSA_RX:VSSA_TX:VSS 0.115763f
c_5225 X290/X12/X50/X5/noxref_5 VSSA_RX:VSSA_TX:VSS 0.115615f
c_5229 X290/X12/X50/X5/noxref_6 VSSA_RX:VSSA_TX:VSS 0.115606f
c_5233 X290/X12/X50/X5/noxref_7 VSSA_RX:VSSA_TX:VSS 0.115594f
c_5236 X290/X12/X50/X5/noxref_8 VSSA_RX:VSSA_TX:VSS 0.115763f
c_5241 XI2/XI0/XOP/N1N21 VSSA_RX:VSSA_TX:VSS 0.044969f
c_5258 XI2/XI0/XOP/N10 VSSA_RX:VSSA_TX:VSS 0.872675f
c_5279 XI2/XI0/XOP/N9 VSSA_RX:VSSA_TX:VSS 0.813483f
c_5284 XI2/XI0/XOP/N1N4 VSSA_RX:VSSA_TX:VSS 0.178495f
c_5289 XI2/XI0/XOP/N1N22 VSSA_RX:VSSA_TX:VSS 0.0280327f
c_5307 XI2/XI0/XOP/N8 VSSA_RX:VSSA_TX:VSS 1.5951f
c_5312 XI2/XI0/XOP/N1N24 VSSA_RX:VSSA_TX:VSS 0.0242151f
c_5325 XI2/XI0/XOP/N7 VSSA_RX:VSSA_TX:VSS 0.979187f
c_5334 XI2/XI0/XOP/N3 VSSA_RX:VSSA_TX:VSS 0.16487f
c_5338 XI2/XI0/XOP/N4 VSSA_RX:VSSA_TX:VSS 0.204557f
c_5350 XI2/XI0/XOP/N1 VSSA_RX:VSSA_TX:VSS 0.231102f
c_5355 XI2/XI0/XOP/N5 VSSA_RX:VSSA_TX:VSS 0.207911f
c_5366 XI2/XI0/XOP/N2 VSSA_RX:VSSA_TX:VSS 0.230379f
c_5370 XI2/XI0/XOP/XI0/N1N5 VSSA_RX:VSSA_TX:VSS 0.0164764f
c_5377 XI2/XI0/XOP/XI0/N4 VSSA_RX:VSSA_TX:VSS 0.151757f
c_5385 XI2/XI0/XOP/XI0/N2 VSSA_RX:VSSA_TX:VSS 0.510439f
c_5391 XI2/XI0/XOP/XI0/N3 VSSA_RX:VSSA_TX:VSS 0.263342f
c_5399 XI2/XI0/XOP/XI0/TIEL VSSA_RX:VSSA_TX:VSS 0.171984f
c_5407 XI2/XI0/XOP/XI0/X1I44/N1N50 VSSA_RX:VSSA_TX:VSS 0.149865f
c_5433 XI2/XI1/TIEH5 VSSA_RX:VSSA_TX:VSS 0.636125f
c_5456 XI2/XI1/TIEH4 VSSA_RX:VSSA_TX:VSS 0.597048f
c_5476 XI2/XI1/TIEH3 VSSA_RX:VSSA_TX:VSS 0.462251f
c_5502 XI2/XI1/TIEH2 VSSA_RX:VSSA_TX:VSS 0.98869f
c_5516 XI2/GMOUT VSSA_RX:VSSA_TX:VSS 22.9815f
c_5525 XI2/XI1/N1N209 VSSA_RX:VSSA_TX:VSS 18.4521f
c_5567 XI2/XI1/VBP VSSA_RX:VSSA_TX:VSS 3.10071f
c_5577 XI2/XI1/N2N77 VSSA_RX:VSSA_TX:VSS 0.375432f
c_5585 XI2/XI1/N2 VSSA_RX:VSSA_TX:VSS 0.556517f
c_5591 XI2/XI1/PDB VSSA_RX:VSSA_TX:VSS 0.10016f
c_5607 XI2/XI1/TIEH1 VSSA_RX:VSSA_TX:VSS 0.306911f
c_5648 XI2/XI1/PDTXB VSSA_RX:VSSA_TX:VSS 2.50463f
c_5662 XI2/XI1/N2N4 VSSA_RX:VSSA_TX:VSS 0.499223f
c_5675 XI2/XI1/X1I241/N1N42 VSSA_RX:VSSA_TX:VSS 0.140075f
c_5678 X290/X13/X6/noxref_30 VSSA_RX:VSSA_TX:VSS 0.0206478f
c_5685 XI2/XI1/N1 VSSA_RX:VSSA_TX:VSS 0.272903f
c_5693 XI2/XI1/N2N116 VSSA_RX:VSSA_TX:VSS 0.204117f
c_5707 XI2/XI1/N2N5 VSSA_RX:VSSA_TX:VSS 0.406933f
c_5716 XI2/XI1/S0B VSSA_RX:VSSA_TX:VSS 0.450924f
c_5726 XI2/XI1/S0 VSSA_RX:VSSA_TX:VSS 0.610105f
c_5731 XI2/XI1/XG9/N1 VSSA_RX:VSSA_TX:VSS 3.18357e-19
c_5745 XI2/XI1/N2N42 VSSA_RX:VSSA_TX:VSS 0.66314f
c_5758 XI2/XI1/N2N95 VSSA_RX:VSSA_TX:VSS 0.188947f
c_5772 XI2/XI1/S2B VSSA_RX:VSSA_TX:VSS 0.417438f
c_5787 XI2/XI1/S2 VSSA_RX:VSSA_TX:VSS 0.563981f
c_5792 XI2/XI1/XG3/N1 VSSA_RX:VSSA_TX:VSS 5.30285e-19
c_5803 XI2/XI1/N1N83 VSSA_RX:VSSA_TX:VSS 0.540507f
c_5811 XI2/XI1/PDRXB VSSA_RX:VSSA_TX:VSS 0.14315f
c_5823 XI2/XI1/N2N69 VSSA_RX:VSSA_TX:VSS 0.460332f
c_5834 XI2/XI1/N2N102 VSSA_RX:VSSA_TX:VSS 0.190054f
c_5846 XI2/XI1/S1B VSSA_RX:VSSA_TX:VSS 0.42132f
c_5859 XI2/XI1/S1 VSSA_RX:VSSA_TX:VSS 0.569586f
c_5864 XI2/XI1/XG6/N1 VSSA_RX:VSSA_TX:VSS 6.08938e-19
c_5868 X290/X13/X7/noxref_6 VSSA_RX:VSSA_TX:VSS 0.11322f
c_5872 X290/X13/X7/noxref_7 VSSA_RX:VSSA_TX:VSS 0.111064f
c_5876 X290/X13/X7/noxref_8 VSSA_RX:VSSA_TX:VSS 0.113105f
c_5880 X290/X13/X7/noxref_9 VSSA_RX:VSSA_TX:VSS 0.111064f
c_5884 X290/X13/X7/noxref_10 VSSA_RX:VSSA_TX:VSS 0.113105f
c_5888 X290/X13/X7/noxref_11 VSSA_RX:VSSA_TX:VSS 0.111064f
c_5892 X290/X13/X7/noxref_12 VSSA_RX:VSSA_TX:VSS 0.113105f
c_5895 X290/X13/X7/noxref_13 VSSA_RX:VSSA_TX:VSS 0.111064f
c_5899 X290/X13/X7/noxref_14 VSSA_RX:VSSA_TX:VSS 0.113212f
c_5913 XI2/XI1/X2I178/N1N42 VSSA_RX:VSSA_TX:VSS 0.252574f
c_5927 XI2/XI1/X2I176/N1N42 VSSA_RX:VSSA_TX:VSS 0.213847f
c_5940 XI2/XI1/X2I174/N1N42 VSSA_RX:VSSA_TX:VSS 0.207617f
c_5951 XI2/XI1/X2I171/N1N42 VSSA_RX:VSSA_TX:VSS 0.251693f
*
.include 'X122G001C_CCW.pex.netlist.X122G001C.pxi'
*
.ends
*
*
